module DivSqrtRecF64_mulAddZ31
(
  clk,
  reset,
  io_inReady_div,
  io_inReady_sqrt,
  io_inValid,
  io_sqrtOp,
  io_a,
  io_b,
  io_roundingMode,
  io_outValid_div,
  io_outValid_sqrt,
  io_out,
  io_exceptionFlags,
  io_usingMulAdd,
  io_latchMulAddA_0,
  io_mulAddA_0,
  io_latchMulAddB_0,
  io_mulAddB_0,
  io_mulAddC_2,
  io_mulAddResult_3
);

  input [64:0] io_a;
  input [64:0] io_b;
  input [1:0] io_roundingMode;
  output [64:0] io_out;
  output [4:0] io_exceptionFlags;
  output [3:0] io_usingMulAdd;
  output [53:0] io_mulAddA_0;
  output [53:0] io_mulAddB_0;
  output [104:0] io_mulAddC_2;
  input [104:0] io_mulAddResult_3;
  input clk;
  input reset;
  input io_inValid;
  input io_sqrtOp;
  output io_inReady_div;
  output io_inReady_sqrt;
  output io_outValid_div;
  output io_outValid_sqrt;
  output io_latchMulAddA_0;
  output io_latchMulAddB_0;
  wire [64:0] io_out;
  wire [4:0] io_exceptionFlags;
  wire [3:0] io_usingMulAdd,T76,T77,T586;
  wire [53:0] io_mulAddA_0,io_mulAddB_0,sigT_C1,zComplSigT_C1,T162,T163,zComplSigT_C1_sqrt,
  T485,T703,sigAdjT_E,T728;
  wire [104:0] io_mulAddC_2,T204,T216,T228;
  wire io_inReady_div,io_inReady_sqrt,io_outValid_div,io_outValid_sqrt,
  io_latchMulAddA_0,io_latchMulAddB_0,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,cyc_E3_sqrt,N119,T13,N120,cyc_C1_div,E_C1_div,T15,
  entering_PC,T17,N121,entering_PB,T19,N122,entering_PA,entering_PA_normalCase,T21,
  cyc_S,T22,T23,ready_PB,T122,valid_leaving_PB,normalCase_PB,N123,ready_PC,T65,
  valid_leaving_PC,T32,T30,normalCase_PC,N124,T54,T33,T40,T34,T49,T41,T47,T48,T52,T50,
  T62,T55,T57,sign_S,T58,T60,T64,T63,T67,leaving_PC,T106,N125,T104,N126,T102,T83,
  N127,cyc_A7_sqrt,cyc_S_sqrt,normalCase_S_sqrt,T87,T86,T89,T88,T91,cyc_S_div,
  normalCase_S_div,T94,T93,T96,T95,T98,T97,T101,T100,T117,T108,T110,T109,T112,T111,T115,
  T113,T119,T118,T121,T120,T124,leaving_PA,valid_leaving_PA,normalCase_PA,N128,
  valid_normalCase_leaving_PA,cyc_B4_div,T129,T128,T140,T131,T133,T132,T135,T134,T138,
  T136,T142,T141,T144,T143,entering_PB_S,T150,T145,leaving_PB,T146,T148,T147,T152,
  T151,T153,normalCase_S,T155,entering_PC_S,T156,T158,T157,T160,T159,T161,T165,
  N129,T166,cyc_C1_sqrt,T167,N130,entering_PC_normalCase,entering_PB_normalCase,T177,
  T178,T180,T183,N131,T198_13,T212,N132,cyc_E3_div,T213,T215,T225,N133,T221,T222,
  cyc_C3_sqrt,cyc_C5_div,T223,cyc_C4_sqrt,cyc_B6_sqrt,N134,cyc_A1_sqrt,N135,
  cyc_A1_div,N136,T269,T262,N137,T267,N138,T270,N139,T281,N140,T280,cyc_A3_sqrt,T287,N141,
  T289,cyc_A3_div,T288,T297,T298,T305_0,zLinPiece_7_A4_div,zLinPiece_6_A4_div,
  zLinPiece_5_A4_div,zLinPiece_4_A4_div,zLinPiece_3_A4_div,zLinPiece_2_A4_div,
  zLinPiece_1_A4_div,zLinPiece_0_A4_div,T339_0,zQuadPiece_3_A6_sqrt,T344,
  zQuadPiece_2_A6_sqrt,T350,T348,zQuadPiece_1_A6_sqrt,T355,T356,zQuadPiece_0_A6_sqrt,T361,T359,
  T362,zQuadPiece_3_A7_sqrt,T367,zQuadPiece_2_A7_sqrt,T373,T371,zQuadPiece_1_A7_sqrt,
  T378,T379,zQuadPiece_0_A7_sqrt,T384,T382,T385,T407,N142,T403,N143,T404,T405,
  cyc_A4,T406,T450,N144,T445,N145,T430,N146,T435,N147,N148,T446,T447,T448,T449,N149,
  T468,T478,T479,T480,T481,T482,N150,N151,N152,cyc_C5_sqrt,cyc_C4_div,N153,T498,T502,
  N154,cyc_B6_div,N155,T512,T511,T515,N156,T519,T520,T521,T522,T523,T524,T530,
  cyc_B2_sqrt,T532,T533,T535,cyc_B1_sqrt,T537,cyc_B3_sqrt,T538,T540,T541,T542,T545,
  T546,T549,cyc_B1_div,T548,T550,T553,cyc_B4_sqrt,T552,T554,T555,T556,T558,
  cyc_A2_div,T559,T561,T562,T565,cyc_B2_div,T564,T566,T569,cyc_B5_sqrt,T568,T570,T571,T572,
  T574,T575,T705,T579,inexactY_E1,hiRoundPosBit_E1,anyRoundExtra_E1,T676,T580,T601,
  N157,T603,T602,T605,N158,T606,T618_13,T618_11,T618_9,T618_7,T618_5,T618_3,
  T618_1,T619_12,T619_10,T619_8,T619_6,T619_4,T619_2,T622_11,T622_10,T622_7,T622_6,
  T622_3,T622_2,T623_9,T623_8,T623_5,T623_4,T626_7,T626_6,T626_5,T626_4,T643_29,
  T643_27,T643_25,T643_23,T643_21,T643_19,T643_17,T643_15,T643_13,T643_11,T643_9,T643_7,
  T643_5,T643_3,T643_1,T644_28,T644_26,T644_24,T644_22,T644_20,T644_18,T644_16,
  T644_14,T644_12,T644_10,T644_8,T644_6,T644_4,T644_2,T647_27,T647_26,T647_23,T647_22,
  T647_19,T647_18,T647_15,T647_14,T647_11,T647_10,T647_7,T647_6,T647_3,T647_2,
  T648_25,T648_24,T648_21,T648_20,T648_17,T648_16,T648_13,T648_12,T648_9,T648_8,
  T648_5,T648_4,T651_23,T651_22,T651_21,T651_20,T651_15,T651_14,T651_13,T651_12,T651_7,
  T651_6,T651_5,T651_4,T652_19,T652_18,T652_17,T652_16,T652_11,T652_10,T652_9,
  T652_8,T655_15,T655_14,T655_13,T655_12,T655_11,T655_10,T655_9,T655_8,T678,T677,T680,
  T681,T684,T688,T689,T690,T691,trueLtX_E1,T696,T693,T698,T697,underflowY_E1,
  totalUnderflowY_E1,T706,T707,T708,T713,N159,sigY_E1_53,T724_53,T715_53,
  roundEvenMask_E1_53,T716,N160,T718,T717,T730,N161,sigY1_E_53,sigY0_E_53,N162,T742,T731,T732,
  T736,T733,T734,T735,T737,T740,T738,T741,T753,T743,T744,T749,T745,all1sHiRoundT_E,
  T746,T747,T751,T750,T752,T754,T756,T755,roundMagDown_PC,T758,T757,T761,N163,T763,
  T762,T764,T768,N164,T769,T770,T773,N165,overflowY_E1,T778,T776,T781,T783,T782,
  T785,T784,T798,notSigNaN_invalid_PC,T793,T786,T792,T787,isInfA_PC,isInfB_PC,T788,
  T790,T794,T796,T795,isNaNB_PC,T800,isSigNaNB_PC,T799,T809,isSigNaNA_PC,isNaNA_PC,
  T801,T803,T806,T813,T814,T815,T817_0,T818,overflowY_roundMagUp_PC,T820,N166,T821,
  notSpecial_isZeroOut_E1,T822,T825,T823,T824,notNaN_isInfOut_E1,T829,T831,T830,
  pegMinFiniteMagOut_E1,T836,T851,T849,T850,T854,T857,T856,T859,T858,T861,T860,T863,
  T862,ready_PA,T864,T866,T869,T868,T871,T870,T873,T872,T875,T874,T877,T876,T879,
  T878,T881,T880,T883,T882,T884,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,
  SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,
  SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,
  SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11,
  SV2V_UNCONNECTED_12,SV2V_UNCONNECTED_13,SV2V_UNCONNECTED_14,
  SV2V_UNCONNECTED_15,SV2V_UNCONNECTED_16,SV2V_UNCONNECTED_17,
  SV2V_UNCONNECTED_18,SV2V_UNCONNECTED_19,SV2V_UNCONNECTED_20,SV2V_UNCONNECTED_21,
  SV2V_UNCONNECTED_22,SV2V_UNCONNECTED_23,SV2V_UNCONNECTED_24,
  SV2V_UNCONNECTED_25,SV2V_UNCONNECTED_26,SV2V_UNCONNECTED_27,
  SV2V_UNCONNECTED_28,SV2V_UNCONNECTED_29,SV2V_UNCONNECTED_30,SV2V_UNCONNECTED_31,
  SV2V_UNCONNECTED_32,SV2V_UNCONNECTED_33,SV2V_UNCONNECTED_34,
  SV2V_UNCONNECTED_35,SV2V_UNCONNECTED_36,SV2V_UNCONNECTED_37,
  SV2V_UNCONNECTED_38,SV2V_UNCONNECTED_39,SV2V_UNCONNECTED_40,SV2V_UNCONNECTED_41,
  SV2V_UNCONNECTED_42,SV2V_UNCONNECTED_43,SV2V_UNCONNECTED_44,
  SV2V_UNCONNECTED_45,SV2V_UNCONNECTED_46,SV2V_UNCONNECTED_47,
  SV2V_UNCONNECTED_48,SV2V_UNCONNECTED_49,SV2V_UNCONNECTED_50,SV2V_UNCONNECTED_51,
  SV2V_UNCONNECTED_52,SV2V_UNCONNECTED_53,SV2V_UNCONNECTED_54,
  SV2V_UNCONNECTED_55,SV2V_UNCONNECTED_56,SV2V_UNCONNECTED_57,
  SV2V_UNCONNECTED_58,SV2V_UNCONNECTED_59,SV2V_UNCONNECTED_60,SV2V_UNCONNECTED_61,
  SV2V_UNCONNECTED_62,SV2V_UNCONNECTED_63,SV2V_UNCONNECTED_64,
  SV2V_UNCONNECTED_65,SV2V_UNCONNECTED_66,SV2V_UNCONNECTED_67,
  SV2V_UNCONNECTED_68,SV2V_UNCONNECTED_69,SV2V_UNCONNECTED_70,SV2V_UNCONNECTED_71,
  SV2V_UNCONNECTED_72,SV2V_UNCONNECTED_73,SV2V_UNCONNECTED_74,
  SV2V_UNCONNECTED_75,SV2V_UNCONNECTED_76,SV2V_UNCONNECTED_77,
  SV2V_UNCONNECTED_78,SV2V_UNCONNECTED_79,SV2V_UNCONNECTED_80,SV2V_UNCONNECTED_81,
  SV2V_UNCONNECTED_82,SV2V_UNCONNECTED_83,SV2V_UNCONNECTED_84,
  SV2V_UNCONNECTED_85,SV2V_UNCONNECTED_86,SV2V_UNCONNECTED_87,
  SV2V_UNCONNECTED_88,SV2V_UNCONNECTED_89,SV2V_UNCONNECTED_90,SV2V_UNCONNECTED_91,
  SV2V_UNCONNECTED_92,SV2V_UNCONNECTED_93,SV2V_UNCONNECTED_94,
  SV2V_UNCONNECTED_95,SV2V_UNCONNECTED_96,SV2V_UNCONNECTED_97,
  SV2V_UNCONNECTED_98,SV2V_UNCONNECTED_99,SV2V_UNCONNECTED_100,SV2V_UNCONNECTED_101,
  SV2V_UNCONNECTED_102,SV2V_UNCONNECTED_103,SV2V_UNCONNECTED_104,
  SV2V_UNCONNECTED_105,SV2V_UNCONNECTED_106,SV2V_UNCONNECTED_107,
  SV2V_UNCONNECTED_108,SV2V_UNCONNECTED_109,SV2V_UNCONNECTED_110,
  SV2V_UNCONNECTED_111,SV2V_UNCONNECTED_112,SV2V_UNCONNECTED_113,
  SV2V_UNCONNECTED_114,SV2V_UNCONNECTED_115,SV2V_UNCONNECTED_116,SV2V_UNCONNECTED_117,
  SV2V_UNCONNECTED_118,SV2V_UNCONNECTED_119,SV2V_UNCONNECTED_120,
  SV2V_UNCONNECTED_121,SV2V_UNCONNECTED_122,SV2V_UNCONNECTED_123,
  SV2V_UNCONNECTED_124,SV2V_UNCONNECTED_125,SV2V_UNCONNECTED_126,
  SV2V_UNCONNECTED_127,SV2V_UNCONNECTED_128,SV2V_UNCONNECTED_129,
  SV2V_UNCONNECTED_130,SV2V_UNCONNECTED_131,SV2V_UNCONNECTED_132,SV2V_UNCONNECTED_133,
  SV2V_UNCONNECTED_134,SV2V_UNCONNECTED_135,SV2V_UNCONNECTED_136,
  SV2V_UNCONNECTED_137,SV2V_UNCONNECTED_138,SV2V_UNCONNECTED_139,
  SV2V_UNCONNECTED_140,SV2V_UNCONNECTED_141,SV2V_UNCONNECTED_142,
  SV2V_UNCONNECTED_143,SV2V_UNCONNECTED_144,SV2V_UNCONNECTED_145,
  SV2V_UNCONNECTED_146,SV2V_UNCONNECTED_147,SV2V_UNCONNECTED_148,SV2V_UNCONNECTED_149,
  SV2V_UNCONNECTED_150,SV2V_UNCONNECTED_151,SV2V_UNCONNECTED_152,
  SV2V_UNCONNECTED_153,SV2V_UNCONNECTED_154,SV2V_UNCONNECTED_155,
  SV2V_UNCONNECTED_156,SV2V_UNCONNECTED_157,SV2V_UNCONNECTED_158,
  SV2V_UNCONNECTED_159,SV2V_UNCONNECTED_160,SV2V_UNCONNECTED_161,
  SV2V_UNCONNECTED_162,SV2V_UNCONNECTED_163,SV2V_UNCONNECTED_164,SV2V_UNCONNECTED_165,
  SV2V_UNCONNECTED_166,SV2V_UNCONNECTED_167,SV2V_UNCONNECTED_168,
  SV2V_UNCONNECTED_169,SV2V_UNCONNECTED_170,SV2V_UNCONNECTED_171,
  SV2V_UNCONNECTED_172,SV2V_UNCONNECTED_173,SV2V_UNCONNECTED_174,
  SV2V_UNCONNECTED_175,SV2V_UNCONNECTED_176,SV2V_UNCONNECTED_177,
  SV2V_UNCONNECTED_178,SV2V_UNCONNECTED_179,SV2V_UNCONNECTED_180,SV2V_UNCONNECTED_181,
  SV2V_UNCONNECTED_182,SV2V_UNCONNECTED_183,SV2V_UNCONNECTED_184,
  SV2V_UNCONNECTED_185,SV2V_UNCONNECTED_186,SV2V_UNCONNECTED_187,
  SV2V_UNCONNECTED_188,SV2V_UNCONNECTED_189,SV2V_UNCONNECTED_190,
  SV2V_UNCONNECTED_191,SV2V_UNCONNECTED_192,SV2V_UNCONNECTED_193,
  SV2V_UNCONNECTED_194,SV2V_UNCONNECTED_195,SV2V_UNCONNECTED_196,SV2V_UNCONNECTED_197,
  SV2V_UNCONNECTED_198,SV2V_UNCONNECTED_199,SV2V_UNCONNECTED_200,
  SV2V_UNCONNECTED_201,SV2V_UNCONNECTED_202,SV2V_UNCONNECTED_203,
  SV2V_UNCONNECTED_204,SV2V_UNCONNECTED_205,SV2V_UNCONNECTED_206,
  SV2V_UNCONNECTED_207,SV2V_UNCONNECTED_208,SV2V_UNCONNECTED_209,
  SV2V_UNCONNECTED_210,SV2V_UNCONNECTED_211,SV2V_UNCONNECTED_212,SV2V_UNCONNECTED_213,
  SV2V_UNCONNECTED_214,SV2V_UNCONNECTED_215,SV2V_UNCONNECTED_216,
  SV2V_UNCONNECTED_217,SV2V_UNCONNECTED_218,SV2V_UNCONNECTED_219,
  SV2V_UNCONNECTED_220,SV2V_UNCONNECTED_221,SV2V_UNCONNECTED_222,
  SV2V_UNCONNECTED_223,SV2V_UNCONNECTED_224,SV2V_UNCONNECTED_225,
  SV2V_UNCONNECTED_226,SV2V_UNCONNECTED_227,SV2V_UNCONNECTED_228,SV2V_UNCONNECTED_229,
  SV2V_UNCONNECTED_230,SV2V_UNCONNECTED_231,SV2V_UNCONNECTED_232,
  SV2V_UNCONNECTED_233,SV2V_UNCONNECTED_234,SV2V_UNCONNECTED_235,
  SV2V_UNCONNECTED_236,SV2V_UNCONNECTED_237,SV2V_UNCONNECTED_238,
  SV2V_UNCONNECTED_239,SV2V_UNCONNECTED_240,SV2V_UNCONNECTED_241,
  SV2V_UNCONNECTED_242,SV2V_UNCONNECTED_243,SV2V_UNCONNECTED_244,SV2V_UNCONNECTED_245,
  SV2V_UNCONNECTED_246,SV2V_UNCONNECTED_247,SV2V_UNCONNECTED_248,
  SV2V_UNCONNECTED_249,SV2V_UNCONNECTED_250,SV2V_UNCONNECTED_251,
  SV2V_UNCONNECTED_252,SV2V_UNCONNECTED_253,SV2V_UNCONNECTED_254,
  SV2V_UNCONNECTED_255,SV2V_UNCONNECTED_256,SV2V_UNCONNECTED_257,
  SV2V_UNCONNECTED_258,SV2V_UNCONNECTED_259,SV2V_UNCONNECTED_260,SV2V_UNCONNECTED_261,
  SV2V_UNCONNECTED_262,SV2V_UNCONNECTED_263,SV2V_UNCONNECTED_264,
  SV2V_UNCONNECTED_265,SV2V_UNCONNECTED_266,SV2V_UNCONNECTED_267,
  SV2V_UNCONNECTED_268,SV2V_UNCONNECTED_269,SV2V_UNCONNECTED_270,
  SV2V_UNCONNECTED_271,SV2V_UNCONNECTED_272,SV2V_UNCONNECTED_273,
  SV2V_UNCONNECTED_274,SV2V_UNCONNECTED_275,SV2V_UNCONNECTED_276,SV2V_UNCONNECTED_277,
  SV2V_UNCONNECTED_278,SV2V_UNCONNECTED_279,SV2V_UNCONNECTED_280,
  SV2V_UNCONNECTED_281,SV2V_UNCONNECTED_282,SV2V_UNCONNECTED_283,
  SV2V_UNCONNECTED_284,SV2V_UNCONNECTED_285,SV2V_UNCONNECTED_286,
  SV2V_UNCONNECTED_287,SV2V_UNCONNECTED_288,SV2V_UNCONNECTED_289,
  SV2V_UNCONNECTED_290,SV2V_UNCONNECTED_291,SV2V_UNCONNECTED_292,SV2V_UNCONNECTED_293,
  SV2V_UNCONNECTED_294,SV2V_UNCONNECTED_295,SV2V_UNCONNECTED_296,
  SV2V_UNCONNECTED_297,SV2V_UNCONNECTED_298,SV2V_UNCONNECTED_299,
  SV2V_UNCONNECTED_300,SV2V_UNCONNECTED_301,SV2V_UNCONNECTED_302,
  SV2V_UNCONNECTED_303,SV2V_UNCONNECTED_304,SV2V_UNCONNECTED_305,
  SV2V_UNCONNECTED_306,SV2V_UNCONNECTED_307,SV2V_UNCONNECTED_308,SV2V_UNCONNECTED_309,
  SV2V_UNCONNECTED_310,SV2V_UNCONNECTED_311,SV2V_UNCONNECTED_312,
  SV2V_UNCONNECTED_313,SV2V_UNCONNECTED_314,SV2V_UNCONNECTED_315,
  SV2V_UNCONNECTED_316,SV2V_UNCONNECTED_317,SV2V_UNCONNECTED_318,
  SV2V_UNCONNECTED_319,SV2V_UNCONNECTED_320,SV2V_UNCONNECTED_321,
  SV2V_UNCONNECTED_322,SV2V_UNCONNECTED_323,SV2V_UNCONNECTED_324,SV2V_UNCONNECTED_325,
  SV2V_UNCONNECTED_326,SV2V_UNCONNECTED_327,SV2V_UNCONNECTED_328,
  SV2V_UNCONNECTED_329,SV2V_UNCONNECTED_330,SV2V_UNCONNECTED_331,
  SV2V_UNCONNECTED_332,SV2V_UNCONNECTED_333,SV2V_UNCONNECTED_334,
  SV2V_UNCONNECTED_335,SV2V_UNCONNECTED_336,SV2V_UNCONNECTED_337,
  SV2V_UNCONNECTED_338,SV2V_UNCONNECTED_339,SV2V_UNCONNECTED_340,SV2V_UNCONNECTED_341,
  SV2V_UNCONNECTED_342,SV2V_UNCONNECTED_343,SV2V_UNCONNECTED_344,
  SV2V_UNCONNECTED_345,SV2V_UNCONNECTED_346,SV2V_UNCONNECTED_347,
  SV2V_UNCONNECTED_348,SV2V_UNCONNECTED_349,SV2V_UNCONNECTED_350,
  SV2V_UNCONNECTED_351,SV2V_UNCONNECTED_352,SV2V_UNCONNECTED_353,
  SV2V_UNCONNECTED_354,SV2V_UNCONNECTED_355,SV2V_UNCONNECTED_356,SV2V_UNCONNECTED_357,
  SV2V_UNCONNECTED_358,SV2V_UNCONNECTED_359,SV2V_UNCONNECTED_360,
  SV2V_UNCONNECTED_361,SV2V_UNCONNECTED_362,SV2V_UNCONNECTED_363,
  SV2V_UNCONNECTED_364,SV2V_UNCONNECTED_365,SV2V_UNCONNECTED_366,
  SV2V_UNCONNECTED_367,SV2V_UNCONNECTED_368,SV2V_UNCONNECTED_369,
  SV2V_UNCONNECTED_370,SV2V_UNCONNECTED_371,SV2V_UNCONNECTED_372,SV2V_UNCONNECTED_373,
  SV2V_UNCONNECTED_374,SV2V_UNCONNECTED_375,SV2V_UNCONNECTED_376,
  SV2V_UNCONNECTED_377,SV2V_UNCONNECTED_378,SV2V_UNCONNECTED_379,
  SV2V_UNCONNECTED_380,SV2V_UNCONNECTED_381,SV2V_UNCONNECTED_382,
  SV2V_UNCONNECTED_383,SV2V_UNCONNECTED_384,SV2V_UNCONNECTED_385,
  SV2V_UNCONNECTED_386,SV2V_UNCONNECTED_387,SV2V_UNCONNECTED_388,SV2V_UNCONNECTED_389,
  SV2V_UNCONNECTED_390,SV2V_UNCONNECTED_391,SV2V_UNCONNECTED_392,
  SV2V_UNCONNECTED_393,SV2V_UNCONNECTED_394,SV2V_UNCONNECTED_395,
  SV2V_UNCONNECTED_396,SV2V_UNCONNECTED_397,SV2V_UNCONNECTED_398,
  SV2V_UNCONNECTED_399,SV2V_UNCONNECTED_400,SV2V_UNCONNECTED_401,
  SV2V_UNCONNECTED_402,SV2V_UNCONNECTED_403,SV2V_UNCONNECTED_404,SV2V_UNCONNECTED_405,
  SV2V_UNCONNECTED_406,SV2V_UNCONNECTED_407,SV2V_UNCONNECTED_408,
  SV2V_UNCONNECTED_409,SV2V_UNCONNECTED_410,SV2V_UNCONNECTED_411,
  SV2V_UNCONNECTED_412,SV2V_UNCONNECTED_413,SV2V_UNCONNECTED_414,
  SV2V_UNCONNECTED_415,SV2V_UNCONNECTED_416,SV2V_UNCONNECTED_417,
  SV2V_UNCONNECTED_418,SV2V_UNCONNECTED_419,SV2V_UNCONNECTED_420,SV2V_UNCONNECTED_421,
  SV2V_UNCONNECTED_422,SV2V_UNCONNECTED_423,SV2V_UNCONNECTED_424,
  SV2V_UNCONNECTED_425,SV2V_UNCONNECTED_426,SV2V_UNCONNECTED_427,
  SV2V_UNCONNECTED_428,SV2V_UNCONNECTED_429,SV2V_UNCONNECTED_430,
  SV2V_UNCONNECTED_431,SV2V_UNCONNECTED_432,SV2V_UNCONNECTED_433,
  SV2V_UNCONNECTED_434,SV2V_UNCONNECTED_435,SV2V_UNCONNECTED_436,SV2V_UNCONNECTED_437,
  SV2V_UNCONNECTED_438,SV2V_UNCONNECTED_439,SV2V_UNCONNECTED_440,
  SV2V_UNCONNECTED_441,SV2V_UNCONNECTED_442,SV2V_UNCONNECTED_443,
  SV2V_UNCONNECTED_444,SV2V_UNCONNECTED_445,SV2V_UNCONNECTED_446,
  SV2V_UNCONNECTED_447,SV2V_UNCONNECTED_448,SV2V_UNCONNECTED_449,
  SV2V_UNCONNECTED_450,SV2V_UNCONNECTED_451,SV2V_UNCONNECTED_452,SV2V_UNCONNECTED_453,
  SV2V_UNCONNECTED_454,SV2V_UNCONNECTED_455,SV2V_UNCONNECTED_456,
  SV2V_UNCONNECTED_457,SV2V_UNCONNECTED_458,SV2V_UNCONNECTED_459,
  SV2V_UNCONNECTED_460,SV2V_UNCONNECTED_461,SV2V_UNCONNECTED_462,
  SV2V_UNCONNECTED_463,SV2V_UNCONNECTED_464,SV2V_UNCONNECTED_465,
  SV2V_UNCONNECTED_466,SV2V_UNCONNECTED_467,SV2V_UNCONNECTED_468,SV2V_UNCONNECTED_469,
  SV2V_UNCONNECTED_470,SV2V_UNCONNECTED_471,SV2V_UNCONNECTED_472,
  SV2V_UNCONNECTED_473,SV2V_UNCONNECTED_474,SV2V_UNCONNECTED_475,
  SV2V_UNCONNECTED_476,SV2V_UNCONNECTED_477,SV2V_UNCONNECTED_478,
  SV2V_UNCONNECTED_479,SV2V_UNCONNECTED_480,SV2V_UNCONNECTED_481,
  SV2V_UNCONNECTED_482,SV2V_UNCONNECTED_483,SV2V_UNCONNECTED_484,SV2V_UNCONNECTED_485,
  SV2V_UNCONNECTED_486,SV2V_UNCONNECTED_487,SV2V_UNCONNECTED_488,
  SV2V_UNCONNECTED_489,SV2V_UNCONNECTED_490,SV2V_UNCONNECTED_491,
  SV2V_UNCONNECTED_492,SV2V_UNCONNECTED_493,SV2V_UNCONNECTED_494,
  SV2V_UNCONNECTED_495,SV2V_UNCONNECTED_496,SV2V_UNCONNECTED_497,
  SV2V_UNCONNECTED_498,SV2V_UNCONNECTED_499,SV2V_UNCONNECTED_500,SV2V_UNCONNECTED_501,
  SV2V_UNCONNECTED_502,SV2V_UNCONNECTED_503,SV2V_UNCONNECTED_504,
  SV2V_UNCONNECTED_505,SV2V_UNCONNECTED_506,SV2V_UNCONNECTED_507,
  SV2V_UNCONNECTED_508,SV2V_UNCONNECTED_509,SV2V_UNCONNECTED_510,
  SV2V_UNCONNECTED_511,SV2V_UNCONNECTED_512,SV2V_UNCONNECTED_513,
  SV2V_UNCONNECTED_514,SV2V_UNCONNECTED_515,SV2V_UNCONNECTED_516,SV2V_UNCONNECTED_517,
  SV2V_UNCONNECTED_518,SV2V_UNCONNECTED_519,SV2V_UNCONNECTED_520,
  SV2V_UNCONNECTED_521,SV2V_UNCONNECTED_522,SV2V_UNCONNECTED_523,
  SV2V_UNCONNECTED_524,SV2V_UNCONNECTED_525,SV2V_UNCONNECTED_526,
  SV2V_UNCONNECTED_527,SV2V_UNCONNECTED_528,SV2V_UNCONNECTED_529,
  SV2V_UNCONNECTED_530,SV2V_UNCONNECTED_531,SV2V_UNCONNECTED_532,SV2V_UNCONNECTED_533,
  SV2V_UNCONNECTED_534,SV2V_UNCONNECTED_535,SV2V_UNCONNECTED_536,
  SV2V_UNCONNECTED_537,SV2V_UNCONNECTED_538,SV2V_UNCONNECTED_539,
  SV2V_UNCONNECTED_540,SV2V_UNCONNECTED_541,SV2V_UNCONNECTED_542,
  SV2V_UNCONNECTED_543,SV2V_UNCONNECTED_544,SV2V_UNCONNECTED_545,
  SV2V_UNCONNECTED_546,SV2V_UNCONNECTED_547,SV2V_UNCONNECTED_548,SV2V_UNCONNECTED_549,
  SV2V_UNCONNECTED_550,SV2V_UNCONNECTED_551,SV2V_UNCONNECTED_552,
  SV2V_UNCONNECTED_553,SV2V_UNCONNECTED_554,SV2V_UNCONNECTED_555,
  SV2V_UNCONNECTED_556,SV2V_UNCONNECTED_557,SV2V_UNCONNECTED_558,
  SV2V_UNCONNECTED_559,SV2V_UNCONNECTED_560,SV2V_UNCONNECTED_561,
  SV2V_UNCONNECTED_562,SV2V_UNCONNECTED_563,SV2V_UNCONNECTED_564,SV2V_UNCONNECTED_565,
  SV2V_UNCONNECTED_566,SV2V_UNCONNECTED_567,SV2V_UNCONNECTED_568,
  SV2V_UNCONNECTED_569,SV2V_UNCONNECTED_570,SV2V_UNCONNECTED_571,
  SV2V_UNCONNECTED_572,SV2V_UNCONNECTED_573,SV2V_UNCONNECTED_574,
  SV2V_UNCONNECTED_575,SV2V_UNCONNECTED_576,SV2V_UNCONNECTED_577,
  SV2V_UNCONNECTED_578,SV2V_UNCONNECTED_579,SV2V_UNCONNECTED_580,SV2V_UNCONNECTED_581,
  SV2V_UNCONNECTED_582,SV2V_UNCONNECTED_583,SV2V_UNCONNECTED_584,
  SV2V_UNCONNECTED_585,SV2V_UNCONNECTED_586,SV2V_UNCONNECTED_587,
  SV2V_UNCONNECTED_588,SV2V_UNCONNECTED_589,SV2V_UNCONNECTED_590,
  SV2V_UNCONNECTED_591,SV2V_UNCONNECTED_592,SV2V_UNCONNECTED_593,
  SV2V_UNCONNECTED_594,SV2V_UNCONNECTED_595,SV2V_UNCONNECTED_596,SV2V_UNCONNECTED_597,
  SV2V_UNCONNECTED_598,SV2V_UNCONNECTED_599,SV2V_UNCONNECTED_600,
  SV2V_UNCONNECTED_601,SV2V_UNCONNECTED_602,SV2V_UNCONNECTED_603,
  SV2V_UNCONNECTED_604,SV2V_UNCONNECTED_605,SV2V_UNCONNECTED_606,
  SV2V_UNCONNECTED_607,SV2V_UNCONNECTED_608,SV2V_UNCONNECTED_609,
  SV2V_UNCONNECTED_610,SV2V_UNCONNECTED_611,SV2V_UNCONNECTED_612,SV2V_UNCONNECTED_613,
  SV2V_UNCONNECTED_614,SV2V_UNCONNECTED_615,SV2V_UNCONNECTED_616,
  SV2V_UNCONNECTED_617,SV2V_UNCONNECTED_618,SV2V_UNCONNECTED_619,
  SV2V_UNCONNECTED_620,SV2V_UNCONNECTED_621,SV2V_UNCONNECTED_622,
  SV2V_UNCONNECTED_623,SV2V_UNCONNECTED_624,SV2V_UNCONNECTED_625,
  SV2V_UNCONNECTED_626,SV2V_UNCONNECTED_627,SV2V_UNCONNECTED_628,SV2V_UNCONNECTED_629,
  SV2V_UNCONNECTED_630,SV2V_UNCONNECTED_631,SV2V_UNCONNECTED_632,
  SV2V_UNCONNECTED_633,SV2V_UNCONNECTED_634,SV2V_UNCONNECTED_635,
  SV2V_UNCONNECTED_636,SV2V_UNCONNECTED_637,SV2V_UNCONNECTED_638,
  SV2V_UNCONNECTED_639,SV2V_UNCONNECTED_640,SV2V_UNCONNECTED_641,
  SV2V_UNCONNECTED_642,SV2V_UNCONNECTED_643,SV2V_UNCONNECTED_644,SV2V_UNCONNECTED_645,
  SV2V_UNCONNECTED_646,SV2V_UNCONNECTED_647,SV2V_UNCONNECTED_648,
  SV2V_UNCONNECTED_649,SV2V_UNCONNECTED_650,SV2V_UNCONNECTED_651,
  SV2V_UNCONNECTED_652,SV2V_UNCONNECTED_653,SV2V_UNCONNECTED_654,
  SV2V_UNCONNECTED_655,SV2V_UNCONNECTED_656,SV2V_UNCONNECTED_657,
  SV2V_UNCONNECTED_658,SV2V_UNCONNECTED_659,SV2V_UNCONNECTED_660,SV2V_UNCONNECTED_661,
  SV2V_UNCONNECTED_662,SV2V_UNCONNECTED_663,SV2V_UNCONNECTED_664,
  SV2V_UNCONNECTED_665,SV2V_UNCONNECTED_666,SV2V_UNCONNECTED_667,
  SV2V_UNCONNECTED_668,SV2V_UNCONNECTED_669,SV2V_UNCONNECTED_670,
  SV2V_UNCONNECTED_671,SV2V_UNCONNECTED_672,SV2V_UNCONNECTED_673,
  SV2V_UNCONNECTED_674,SV2V_UNCONNECTED_675,SV2V_UNCONNECTED_676,SV2V_UNCONNECTED_677,
  SV2V_UNCONNECTED_678,SV2V_UNCONNECTED_679,SV2V_UNCONNECTED_680,
  SV2V_UNCONNECTED_681,SV2V_UNCONNECTED_682,SV2V_UNCONNECTED_683,
  SV2V_UNCONNECTED_684,SV2V_UNCONNECTED_685,SV2V_UNCONNECTED_686,
  SV2V_UNCONNECTED_687,SV2V_UNCONNECTED_688,SV2V_UNCONNECTED_689,
  SV2V_UNCONNECTED_690,SV2V_UNCONNECTED_691,SV2V_UNCONNECTED_692,SV2V_UNCONNECTED_693,
  SV2V_UNCONNECTED_694,SV2V_UNCONNECTED_695,SV2V_UNCONNECTED_696,
  SV2V_UNCONNECTED_697,SV2V_UNCONNECTED_698,SV2V_UNCONNECTED_699,
  SV2V_UNCONNECTED_700,SV2V_UNCONNECTED_701,SV2V_UNCONNECTED_702,
  SV2V_UNCONNECTED_703,SV2V_UNCONNECTED_704,SV2V_UNCONNECTED_705,
  SV2V_UNCONNECTED_706,SV2V_UNCONNECTED_707,SV2V_UNCONNECTED_708,SV2V_UNCONNECTED_709,
  SV2V_UNCONNECTED_710,SV2V_UNCONNECTED_711,SV2V_UNCONNECTED_712,
  SV2V_UNCONNECTED_713,SV2V_UNCONNECTED_714,SV2V_UNCONNECTED_715,
  SV2V_UNCONNECTED_716,SV2V_UNCONNECTED_717,SV2V_UNCONNECTED_718,
  SV2V_UNCONNECTED_719,SV2V_UNCONNECTED_720,SV2V_UNCONNECTED_721,
  SV2V_UNCONNECTED_722,SV2V_UNCONNECTED_723,SV2V_UNCONNECTED_724,SV2V_UNCONNECTED_725,
  SV2V_UNCONNECTED_726,SV2V_UNCONNECTED_727,SV2V_UNCONNECTED_728,
  SV2V_UNCONNECTED_729,SV2V_UNCONNECTED_730,SV2V_UNCONNECTED_731,
  SV2V_UNCONNECTED_732,SV2V_UNCONNECTED_733,SV2V_UNCONNECTED_734,
  SV2V_UNCONNECTED_735,SV2V_UNCONNECTED_736,SV2V_UNCONNECTED_737,
  SV2V_UNCONNECTED_738,SV2V_UNCONNECTED_739,SV2V_UNCONNECTED_740,SV2V_UNCONNECTED_741,
  SV2V_UNCONNECTED_742,SV2V_UNCONNECTED_743,SV2V_UNCONNECTED_744,
  SV2V_UNCONNECTED_745,SV2V_UNCONNECTED_746,SV2V_UNCONNECTED_747,
  SV2V_UNCONNECTED_748,SV2V_UNCONNECTED_749,SV2V_UNCONNECTED_750,
  SV2V_UNCONNECTED_751,SV2V_UNCONNECTED_752,SV2V_UNCONNECTED_753,
  SV2V_UNCONNECTED_754,SV2V_UNCONNECTED_755,SV2V_UNCONNECTED_756,SV2V_UNCONNECTED_757,
  SV2V_UNCONNECTED_758,SV2V_UNCONNECTED_759,SV2V_UNCONNECTED_760,
  SV2V_UNCONNECTED_761,SV2V_UNCONNECTED_762,SV2V_UNCONNECTED_763,
  SV2V_UNCONNECTED_764,SV2V_UNCONNECTED_765,SV2V_UNCONNECTED_766,
  SV2V_UNCONNECTED_767,SV2V_UNCONNECTED_768,SV2V_UNCONNECTED_769,
  SV2V_UNCONNECTED_770,SV2V_UNCONNECTED_771,SV2V_UNCONNECTED_772,SV2V_UNCONNECTED_773,
  SV2V_UNCONNECTED_774,SV2V_UNCONNECTED_775,SV2V_UNCONNECTED_776,
  SV2V_UNCONNECTED_777,SV2V_UNCONNECTED_778,SV2V_UNCONNECTED_779,
  SV2V_UNCONNECTED_780,SV2V_UNCONNECTED_781,SV2V_UNCONNECTED_782,
  SV2V_UNCONNECTED_783,SV2V_UNCONNECTED_784,SV2V_UNCONNECTED_785,
  SV2V_UNCONNECTED_786,SV2V_UNCONNECTED_787,SV2V_UNCONNECTED_788,SV2V_UNCONNECTED_789,
  SV2V_UNCONNECTED_790,SV2V_UNCONNECTED_791,SV2V_UNCONNECTED_792,
  SV2V_UNCONNECTED_793,SV2V_UNCONNECTED_794,SV2V_UNCONNECTED_795,
  SV2V_UNCONNECTED_796,SV2V_UNCONNECTED_797,SV2V_UNCONNECTED_798,
  SV2V_UNCONNECTED_799,SV2V_UNCONNECTED_800,SV2V_UNCONNECTED_801,
  SV2V_UNCONNECTED_802,SV2V_UNCONNECTED_803,SV2V_UNCONNECTED_804,SV2V_UNCONNECTED_805,
  SV2V_UNCONNECTED_806,SV2V_UNCONNECTED_807,SV2V_UNCONNECTED_808,
  SV2V_UNCONNECTED_809,SV2V_UNCONNECTED_810,SV2V_UNCONNECTED_811,
  SV2V_UNCONNECTED_812,SV2V_UNCONNECTED_813,SV2V_UNCONNECTED_814,
  SV2V_UNCONNECTED_815,SV2V_UNCONNECTED_816,SV2V_UNCONNECTED_817,
  SV2V_UNCONNECTED_818,SV2V_UNCONNECTED_819,SV2V_UNCONNECTED_820,SV2V_UNCONNECTED_821,
  SV2V_UNCONNECTED_822,SV2V_UNCONNECTED_823,SV2V_UNCONNECTED_824,
  SV2V_UNCONNECTED_825,SV2V_UNCONNECTED_826,SV2V_UNCONNECTED_827,
  SV2V_UNCONNECTED_828,SV2V_UNCONNECTED_829,SV2V_UNCONNECTED_830,
  SV2V_UNCONNECTED_831,SV2V_UNCONNECTED_832,SV2V_UNCONNECTED_833,
  SV2V_UNCONNECTED_834,SV2V_UNCONNECTED_835,SV2V_UNCONNECTED_836,SV2V_UNCONNECTED_837,
  SV2V_UNCONNECTED_838,SV2V_UNCONNECTED_839,SV2V_UNCONNECTED_840,
  SV2V_UNCONNECTED_841,SV2V_UNCONNECTED_842,SV2V_UNCONNECTED_843,
  SV2V_UNCONNECTED_844,SV2V_UNCONNECTED_845,SV2V_UNCONNECTED_846,
  SV2V_UNCONNECTED_847,SV2V_UNCONNECTED_848,SV2V_UNCONNECTED_849,
  SV2V_UNCONNECTED_850,SV2V_UNCONNECTED_851,SV2V_UNCONNECTED_852,SV2V_UNCONNECTED_853,
  SV2V_UNCONNECTED_854,SV2V_UNCONNECTED_855,SV2V_UNCONNECTED_856,
  SV2V_UNCONNECTED_857,SV2V_UNCONNECTED_858,SV2V_UNCONNECTED_859,
  SV2V_UNCONNECTED_860,SV2V_UNCONNECTED_861,SV2V_UNCONNECTED_862,
  SV2V_UNCONNECTED_863,SV2V_UNCONNECTED_864,SV2V_UNCONNECTED_865,
  SV2V_UNCONNECTED_866,SV2V_UNCONNECTED_867,SV2V_UNCONNECTED_868,SV2V_UNCONNECTED_869,
  SV2V_UNCONNECTED_870,SV2V_UNCONNECTED_871,SV2V_UNCONNECTED_872,
  SV2V_UNCONNECTED_873,SV2V_UNCONNECTED_874,SV2V_UNCONNECTED_875,
  SV2V_UNCONNECTED_876,SV2V_UNCONNECTED_877,SV2V_UNCONNECTED_878,
  SV2V_UNCONNECTED_879,SV2V_UNCONNECTED_880,SV2V_UNCONNECTED_881,
  SV2V_UNCONNECTED_882,SV2V_UNCONNECTED_883,SV2V_UNCONNECTED_884,SV2V_UNCONNECTED_885,
  SV2V_UNCONNECTED_886,SV2V_UNCONNECTED_887,SV2V_UNCONNECTED_888,
  SV2V_UNCONNECTED_889,SV2V_UNCONNECTED_890,SV2V_UNCONNECTED_891,
  SV2V_UNCONNECTED_892,SV2V_UNCONNECTED_893,SV2V_UNCONNECTED_894,
  SV2V_UNCONNECTED_895,SV2V_UNCONNECTED_896,SV2V_UNCONNECTED_897,
  SV2V_UNCONNECTED_898,SV2V_UNCONNECTED_899,SV2V_UNCONNECTED_900,SV2V_UNCONNECTED_901,
  SV2V_UNCONNECTED_902,SV2V_UNCONNECTED_903,SV2V_UNCONNECTED_904,
  SV2V_UNCONNECTED_905,SV2V_UNCONNECTED_906,SV2V_UNCONNECTED_907,
  SV2V_UNCONNECTED_908,SV2V_UNCONNECTED_909,SV2V_UNCONNECTED_910,
  SV2V_UNCONNECTED_911,SV2V_UNCONNECTED_912,SV2V_UNCONNECTED_913,
  SV2V_UNCONNECTED_914,SV2V_UNCONNECTED_915,SV2V_UNCONNECTED_916,SV2V_UNCONNECTED_917,
  SV2V_UNCONNECTED_918,SV2V_UNCONNECTED_919,SV2V_UNCONNECTED_920,
  SV2V_UNCONNECTED_921,SV2V_UNCONNECTED_922,SV2V_UNCONNECTED_923,
  SV2V_UNCONNECTED_924,SV2V_UNCONNECTED_925,SV2V_UNCONNECTED_926,
  SV2V_UNCONNECTED_927,SV2V_UNCONNECTED_928,SV2V_UNCONNECTED_929,
  SV2V_UNCONNECTED_930,SV2V_UNCONNECTED_931,SV2V_UNCONNECTED_932,SV2V_UNCONNECTED_933,
  SV2V_UNCONNECTED_934,SV2V_UNCONNECTED_935,SV2V_UNCONNECTED_936,
  SV2V_UNCONNECTED_937,SV2V_UNCONNECTED_938,SV2V_UNCONNECTED_939,
  SV2V_UNCONNECTED_940,SV2V_UNCONNECTED_941,SV2V_UNCONNECTED_942,
  SV2V_UNCONNECTED_943,SV2V_UNCONNECTED_944,SV2V_UNCONNECTED_945,
  SV2V_UNCONNECTED_946,SV2V_UNCONNECTED_947,SV2V_UNCONNECTED_948,SV2V_UNCONNECTED_949,
  SV2V_UNCONNECTED_950,SV2V_UNCONNECTED_951,SV2V_UNCONNECTED_952,
  SV2V_UNCONNECTED_953,SV2V_UNCONNECTED_954,SV2V_UNCONNECTED_955,
  SV2V_UNCONNECTED_956,SV2V_UNCONNECTED_957,SV2V_UNCONNECTED_958,
  SV2V_UNCONNECTED_959,SV2V_UNCONNECTED_960,SV2V_UNCONNECTED_961,
  SV2V_UNCONNECTED_962,SV2V_UNCONNECTED_963,SV2V_UNCONNECTED_964,SV2V_UNCONNECTED_965,
  SV2V_UNCONNECTED_966,SV2V_UNCONNECTED_967,SV2V_UNCONNECTED_968,
  SV2V_UNCONNECTED_969,SV2V_UNCONNECTED_970,SV2V_UNCONNECTED_971,
  SV2V_UNCONNECTED_972,SV2V_UNCONNECTED_973,SV2V_UNCONNECTED_974,
  SV2V_UNCONNECTED_975,SV2V_UNCONNECTED_976,SV2V_UNCONNECTED_977,
  SV2V_UNCONNECTED_978,SV2V_UNCONNECTED_979,SV2V_UNCONNECTED_980,SV2V_UNCONNECTED_981,
  SV2V_UNCONNECTED_982,SV2V_UNCONNECTED_983,SV2V_UNCONNECTED_984,
  SV2V_UNCONNECTED_985,SV2V_UNCONNECTED_986,SV2V_UNCONNECTED_987,
  SV2V_UNCONNECTED_988,SV2V_UNCONNECTED_989,SV2V_UNCONNECTED_990,
  SV2V_UNCONNECTED_991,SV2V_UNCONNECTED_992,SV2V_UNCONNECTED_993,
  SV2V_UNCONNECTED_994,SV2V_UNCONNECTED_995,SV2V_UNCONNECTED_996,SV2V_UNCONNECTED_997,
  SV2V_UNCONNECTED_998,SV2V_UNCONNECTED_999,SV2V_UNCONNECTED_1000,
  SV2V_UNCONNECTED_1001,SV2V_UNCONNECTED_1002,SV2V_UNCONNECTED_1003,
  SV2V_UNCONNECTED_1004,SV2V_UNCONNECTED_1005,SV2V_UNCONNECTED_1006,
  SV2V_UNCONNECTED_1007,SV2V_UNCONNECTED_1008,SV2V_UNCONNECTED_1009,
  SV2V_UNCONNECTED_1010,SV2V_UNCONNECTED_1011,SV2V_UNCONNECTED_1012,
  SV2V_UNCONNECTED_1013,SV2V_UNCONNECTED_1014,SV2V_UNCONNECTED_1015,
  SV2V_UNCONNECTED_1016,SV2V_UNCONNECTED_1017,SV2V_UNCONNECTED_1018,
  SV2V_UNCONNECTED_1019,SV2V_UNCONNECTED_1020,SV2V_UNCONNECTED_1021,
  SV2V_UNCONNECTED_1022,SV2V_UNCONNECTED_1023,SV2V_UNCONNECTED_1024,
  SV2V_UNCONNECTED_1025,SV2V_UNCONNECTED_1026,SV2V_UNCONNECTED_1027,SV2V_UNCONNECTED_1028,
  SV2V_UNCONNECTED_1029,SV2V_UNCONNECTED_1030,SV2V_UNCONNECTED_1031,
  SV2V_UNCONNECTED_1032,SV2V_UNCONNECTED_1033,SV2V_UNCONNECTED_1034,
  SV2V_UNCONNECTED_1035,SV2V_UNCONNECTED_1036,SV2V_UNCONNECTED_1037,
  SV2V_UNCONNECTED_1038,SV2V_UNCONNECTED_1039,SV2V_UNCONNECTED_1040,
  SV2V_UNCONNECTED_1041,SV2V_UNCONNECTED_1042,SV2V_UNCONNECTED_1043,
  SV2V_UNCONNECTED_1044,SV2V_UNCONNECTED_1045,SV2V_UNCONNECTED_1046,
  SV2V_UNCONNECTED_1047,SV2V_UNCONNECTED_1048,SV2V_UNCONNECTED_1049,
  SV2V_UNCONNECTED_1050,SV2V_UNCONNECTED_1051,SV2V_UNCONNECTED_1052,
  SV2V_UNCONNECTED_1053,SV2V_UNCONNECTED_1054,SV2V_UNCONNECTED_1055,
  SV2V_UNCONNECTED_1056,SV2V_UNCONNECTED_1057,SV2V_UNCONNECTED_1058,
  SV2V_UNCONNECTED_1059,SV2V_UNCONNECTED_1060,SV2V_UNCONNECTED_1061,
  SV2V_UNCONNECTED_1062,SV2V_UNCONNECTED_1063,SV2V_UNCONNECTED_1064,
  SV2V_UNCONNECTED_1065,SV2V_UNCONNECTED_1066,SV2V_UNCONNECTED_1067,SV2V_UNCONNECTED_1068,
  SV2V_UNCONNECTED_1069,SV2V_UNCONNECTED_1070,SV2V_UNCONNECTED_1071,
  SV2V_UNCONNECTED_1072,SV2V_UNCONNECTED_1073,SV2V_UNCONNECTED_1074,
  SV2V_UNCONNECTED_1075,SV2V_UNCONNECTED_1076,SV2V_UNCONNECTED_1077,
  SV2V_UNCONNECTED_1078,SV2V_UNCONNECTED_1079,SV2V_UNCONNECTED_1080,
  SV2V_UNCONNECTED_1081,SV2V_UNCONNECTED_1082,SV2V_UNCONNECTED_1083,
  SV2V_UNCONNECTED_1084,SV2V_UNCONNECTED_1085,SV2V_UNCONNECTED_1086,
  SV2V_UNCONNECTED_1087,SV2V_UNCONNECTED_1088,SV2V_UNCONNECTED_1089,
  SV2V_UNCONNECTED_1090,SV2V_UNCONNECTED_1091,SV2V_UNCONNECTED_1092,
  SV2V_UNCONNECTED_1093,SV2V_UNCONNECTED_1094,SV2V_UNCONNECTED_1095,
  SV2V_UNCONNECTED_1096,SV2V_UNCONNECTED_1097,SV2V_UNCONNECTED_1098,
  SV2V_UNCONNECTED_1099,SV2V_UNCONNECTED_1100,SV2V_UNCONNECTED_1101,
  SV2V_UNCONNECTED_1102,SV2V_UNCONNECTED_1103,SV2V_UNCONNECTED_1104,
  SV2V_UNCONNECTED_1105,SV2V_UNCONNECTED_1106,SV2V_UNCONNECTED_1107,SV2V_UNCONNECTED_1108,
  SV2V_UNCONNECTED_1109,SV2V_UNCONNECTED_1110,SV2V_UNCONNECTED_1111,
  SV2V_UNCONNECTED_1112,SV2V_UNCONNECTED_1113,SV2V_UNCONNECTED_1114,
  SV2V_UNCONNECTED_1115,SV2V_UNCONNECTED_1116,SV2V_UNCONNECTED_1117,
  SV2V_UNCONNECTED_1118,SV2V_UNCONNECTED_1119,SV2V_UNCONNECTED_1120,
  SV2V_UNCONNECTED_1121,SV2V_UNCONNECTED_1122,SV2V_UNCONNECTED_1123,
  SV2V_UNCONNECTED_1124,SV2V_UNCONNECTED_1125,SV2V_UNCONNECTED_1126,
  SV2V_UNCONNECTED_1127,SV2V_UNCONNECTED_1128,SV2V_UNCONNECTED_1129,
  SV2V_UNCONNECTED_1130,SV2V_UNCONNECTED_1131,SV2V_UNCONNECTED_1132,
  SV2V_UNCONNECTED_1133,SV2V_UNCONNECTED_1134,SV2V_UNCONNECTED_1135,
  SV2V_UNCONNECTED_1136,SV2V_UNCONNECTED_1137,SV2V_UNCONNECTED_1138,
  SV2V_UNCONNECTED_1139,SV2V_UNCONNECTED_1140,SV2V_UNCONNECTED_1141,
  SV2V_UNCONNECTED_1142,SV2V_UNCONNECTED_1143,SV2V_UNCONNECTED_1144,
  SV2V_UNCONNECTED_1145,SV2V_UNCONNECTED_1146,SV2V_UNCONNECTED_1147,SV2V_UNCONNECTED_1148,
  SV2V_UNCONNECTED_1149,SV2V_UNCONNECTED_1150,SV2V_UNCONNECTED_1151,
  SV2V_UNCONNECTED_1152,SV2V_UNCONNECTED_1153,SV2V_UNCONNECTED_1154,
  SV2V_UNCONNECTED_1155,SV2V_UNCONNECTED_1156,SV2V_UNCONNECTED_1157,
  SV2V_UNCONNECTED_1158,SV2V_UNCONNECTED_1159,SV2V_UNCONNECTED_1160,
  SV2V_UNCONNECTED_1161,SV2V_UNCONNECTED_1162,SV2V_UNCONNECTED_1163,
  SV2V_UNCONNECTED_1164,SV2V_UNCONNECTED_1165,SV2V_UNCONNECTED_1166,
  SV2V_UNCONNECTED_1167,SV2V_UNCONNECTED_1168,SV2V_UNCONNECTED_1169,
  SV2V_UNCONNECTED_1170,SV2V_UNCONNECTED_1171,SV2V_UNCONNECTED_1172,
  SV2V_UNCONNECTED_1173,SV2V_UNCONNECTED_1174,SV2V_UNCONNECTED_1175,
  SV2V_UNCONNECTED_1176,SV2V_UNCONNECTED_1177,SV2V_UNCONNECTED_1178,
  SV2V_UNCONNECTED_1179,SV2V_UNCONNECTED_1180,SV2V_UNCONNECTED_1181,
  SV2V_UNCONNECTED_1182,SV2V_UNCONNECTED_1183,SV2V_UNCONNECTED_1184,
  SV2V_UNCONNECTED_1185,SV2V_UNCONNECTED_1186,SV2V_UNCONNECTED_1187,SV2V_UNCONNECTED_1188,
  SV2V_UNCONNECTED_1189,SV2V_UNCONNECTED_1190,SV2V_UNCONNECTED_1191,
  SV2V_UNCONNECTED_1192,SV2V_UNCONNECTED_1193,SV2V_UNCONNECTED_1194,
  SV2V_UNCONNECTED_1195,SV2V_UNCONNECTED_1196,SV2V_UNCONNECTED_1197,
  SV2V_UNCONNECTED_1198,SV2V_UNCONNECTED_1199,SV2V_UNCONNECTED_1200,
  SV2V_UNCONNECTED_1201,SV2V_UNCONNECTED_1202,SV2V_UNCONNECTED_1203,
  SV2V_UNCONNECTED_1204,SV2V_UNCONNECTED_1205,SV2V_UNCONNECTED_1206,
  SV2V_UNCONNECTED_1207,SV2V_UNCONNECTED_1208,SV2V_UNCONNECTED_1209,
  SV2V_UNCONNECTED_1210,SV2V_UNCONNECTED_1211,SV2V_UNCONNECTED_1212,
  SV2V_UNCONNECTED_1213,SV2V_UNCONNECTED_1214,SV2V_UNCONNECTED_1215,
  SV2V_UNCONNECTED_1216,SV2V_UNCONNECTED_1217,SV2V_UNCONNECTED_1218,
  SV2V_UNCONNECTED_1219,SV2V_UNCONNECTED_1220,SV2V_UNCONNECTED_1221,
  SV2V_UNCONNECTED_1222,SV2V_UNCONNECTED_1223,SV2V_UNCONNECTED_1224,
  SV2V_UNCONNECTED_1225,SV2V_UNCONNECTED_1226,SV2V_UNCONNECTED_1227,SV2V_UNCONNECTED_1228,
  SV2V_UNCONNECTED_1229,SV2V_UNCONNECTED_1230,SV2V_UNCONNECTED_1231,
  SV2V_UNCONNECTED_1232,SV2V_UNCONNECTED_1233,SV2V_UNCONNECTED_1234,
  SV2V_UNCONNECTED_1235,SV2V_UNCONNECTED_1236,SV2V_UNCONNECTED_1237,
  SV2V_UNCONNECTED_1238,SV2V_UNCONNECTED_1239,SV2V_UNCONNECTED_1240,
  SV2V_UNCONNECTED_1241,SV2V_UNCONNECTED_1242,SV2V_UNCONNECTED_1243,
  SV2V_UNCONNECTED_1244,SV2V_UNCONNECTED_1245,SV2V_UNCONNECTED_1246,
  SV2V_UNCONNECTED_1247,SV2V_UNCONNECTED_1248,SV2V_UNCONNECTED_1249,
  SV2V_UNCONNECTED_1250,SV2V_UNCONNECTED_1251,SV2V_UNCONNECTED_1252,
  SV2V_UNCONNECTED_1253,SV2V_UNCONNECTED_1254,SV2V_UNCONNECTED_1255,
  SV2V_UNCONNECTED_1256,SV2V_UNCONNECTED_1257,SV2V_UNCONNECTED_1258,
  SV2V_UNCONNECTED_1259,SV2V_UNCONNECTED_1260,SV2V_UNCONNECTED_1261,
  SV2V_UNCONNECTED_1262,SV2V_UNCONNECTED_1263,SV2V_UNCONNECTED_1264,
  SV2V_UNCONNECTED_1265,SV2V_UNCONNECTED_1266,SV2V_UNCONNECTED_1267,SV2V_UNCONNECTED_1268,
  SV2V_UNCONNECTED_1269,SV2V_UNCONNECTED_1270,SV2V_UNCONNECTED_1271,
  SV2V_UNCONNECTED_1272,SV2V_UNCONNECTED_1273,SV2V_UNCONNECTED_1274,
  SV2V_UNCONNECTED_1275,SV2V_UNCONNECTED_1276,SV2V_UNCONNECTED_1277,
  SV2V_UNCONNECTED_1278,SV2V_UNCONNECTED_1279,SV2V_UNCONNECTED_1280,
  SV2V_UNCONNECTED_1281,SV2V_UNCONNECTED_1282,SV2V_UNCONNECTED_1283,
  SV2V_UNCONNECTED_1284,SV2V_UNCONNECTED_1285,SV2V_UNCONNECTED_1286,
  SV2V_UNCONNECTED_1287,SV2V_UNCONNECTED_1288,SV2V_UNCONNECTED_1289,
  SV2V_UNCONNECTED_1290,SV2V_UNCONNECTED_1291,SV2V_UNCONNECTED_1292,
  SV2V_UNCONNECTED_1293,SV2V_UNCONNECTED_1294,SV2V_UNCONNECTED_1295,
  SV2V_UNCONNECTED_1296,SV2V_UNCONNECTED_1297,SV2V_UNCONNECTED_1298,
  SV2V_UNCONNECTED_1299,SV2V_UNCONNECTED_1300,SV2V_UNCONNECTED_1301,
  SV2V_UNCONNECTED_1302,SV2V_UNCONNECTED_1303,SV2V_UNCONNECTED_1304,
  SV2V_UNCONNECTED_1305,SV2V_UNCONNECTED_1306,SV2V_UNCONNECTED_1307,SV2V_UNCONNECTED_1308,
  SV2V_UNCONNECTED_1309,SV2V_UNCONNECTED_1310,SV2V_UNCONNECTED_1311,
  SV2V_UNCONNECTED_1312,SV2V_UNCONNECTED_1313,SV2V_UNCONNECTED_1314,
  SV2V_UNCONNECTED_1315,SV2V_UNCONNECTED_1316,SV2V_UNCONNECTED_1317,
  SV2V_UNCONNECTED_1318,SV2V_UNCONNECTED_1319,SV2V_UNCONNECTED_1320,
  SV2V_UNCONNECTED_1321,SV2V_UNCONNECTED_1322,SV2V_UNCONNECTED_1323,
  SV2V_UNCONNECTED_1324,SV2V_UNCONNECTED_1325,SV2V_UNCONNECTED_1326,
  SV2V_UNCONNECTED_1327,SV2V_UNCONNECTED_1328,SV2V_UNCONNECTED_1329,
  SV2V_UNCONNECTED_1330,SV2V_UNCONNECTED_1331,SV2V_UNCONNECTED_1332,
  SV2V_UNCONNECTED_1333,SV2V_UNCONNECTED_1334,SV2V_UNCONNECTED_1335,
  SV2V_UNCONNECTED_1336,SV2V_UNCONNECTED_1337,SV2V_UNCONNECTED_1338,
  SV2V_UNCONNECTED_1339,SV2V_UNCONNECTED_1340,SV2V_UNCONNECTED_1341,
  SV2V_UNCONNECTED_1342,SV2V_UNCONNECTED_1343,SV2V_UNCONNECTED_1344,
  SV2V_UNCONNECTED_1345,SV2V_UNCONNECTED_1346,SV2V_UNCONNECTED_1347,SV2V_UNCONNECTED_1348,
  SV2V_UNCONNECTED_1349,SV2V_UNCONNECTED_1350,SV2V_UNCONNECTED_1351,
  SV2V_UNCONNECTED_1352,SV2V_UNCONNECTED_1353,SV2V_UNCONNECTED_1354,
  SV2V_UNCONNECTED_1355,SV2V_UNCONNECTED_1356,SV2V_UNCONNECTED_1357,
  SV2V_UNCONNECTED_1358,SV2V_UNCONNECTED_1359,SV2V_UNCONNECTED_1360,
  SV2V_UNCONNECTED_1361,SV2V_UNCONNECTED_1362,SV2V_UNCONNECTED_1363,
  SV2V_UNCONNECTED_1364,SV2V_UNCONNECTED_1365,SV2V_UNCONNECTED_1366,
  SV2V_UNCONNECTED_1367,SV2V_UNCONNECTED_1368,SV2V_UNCONNECTED_1369,
  SV2V_UNCONNECTED_1370,SV2V_UNCONNECTED_1371,SV2V_UNCONNECTED_1372,
  SV2V_UNCONNECTED_1373,SV2V_UNCONNECTED_1374,SV2V_UNCONNECTED_1375,
  SV2V_UNCONNECTED_1376,SV2V_UNCONNECTED_1377,SV2V_UNCONNECTED_1378,
  SV2V_UNCONNECTED_1379,SV2V_UNCONNECTED_1380,SV2V_UNCONNECTED_1381,
  SV2V_UNCONNECTED_1382,SV2V_UNCONNECTED_1383,SV2V_UNCONNECTED_1384,
  SV2V_UNCONNECTED_1385,SV2V_UNCONNECTED_1386,SV2V_UNCONNECTED_1387,SV2V_UNCONNECTED_1388,
  SV2V_UNCONNECTED_1389,SV2V_UNCONNECTED_1390,SV2V_UNCONNECTED_1391,
  SV2V_UNCONNECTED_1392,SV2V_UNCONNECTED_1393,SV2V_UNCONNECTED_1394,
  SV2V_UNCONNECTED_1395,SV2V_UNCONNECTED_1396,SV2V_UNCONNECTED_1397,
  SV2V_UNCONNECTED_1398,SV2V_UNCONNECTED_1399,SV2V_UNCONNECTED_1400,
  SV2V_UNCONNECTED_1401,SV2V_UNCONNECTED_1402,SV2V_UNCONNECTED_1403,
  SV2V_UNCONNECTED_1404,SV2V_UNCONNECTED_1405,SV2V_UNCONNECTED_1406,
  SV2V_UNCONNECTED_1407,SV2V_UNCONNECTED_1408,SV2V_UNCONNECTED_1409,
  SV2V_UNCONNECTED_1410,SV2V_UNCONNECTED_1411,SV2V_UNCONNECTED_1412,
  SV2V_UNCONNECTED_1413,SV2V_UNCONNECTED_1414,SV2V_UNCONNECTED_1415,
  SV2V_UNCONNECTED_1416,SV2V_UNCONNECTED_1417,SV2V_UNCONNECTED_1418,
  SV2V_UNCONNECTED_1419,SV2V_UNCONNECTED_1420,SV2V_UNCONNECTED_1421,
  SV2V_UNCONNECTED_1422,SV2V_UNCONNECTED_1423,SV2V_UNCONNECTED_1424,
  SV2V_UNCONNECTED_1425,SV2V_UNCONNECTED_1426,SV2V_UNCONNECTED_1427,SV2V_UNCONNECTED_1428,
  SV2V_UNCONNECTED_1429,SV2V_UNCONNECTED_1430,SV2V_UNCONNECTED_1431,
  SV2V_UNCONNECTED_1432,SV2V_UNCONNECTED_1433,SV2V_UNCONNECTED_1434,
  SV2V_UNCONNECTED_1435,SV2V_UNCONNECTED_1436,SV2V_UNCONNECTED_1437,
  SV2V_UNCONNECTED_1438,SV2V_UNCONNECTED_1439,SV2V_UNCONNECTED_1440,
  SV2V_UNCONNECTED_1441,SV2V_UNCONNECTED_1442,SV2V_UNCONNECTED_1443,
  SV2V_UNCONNECTED_1444,SV2V_UNCONNECTED_1445,SV2V_UNCONNECTED_1446,
  SV2V_UNCONNECTED_1447,SV2V_UNCONNECTED_1448,SV2V_UNCONNECTED_1449,
  SV2V_UNCONNECTED_1450,SV2V_UNCONNECTED_1451,SV2V_UNCONNECTED_1452,
  SV2V_UNCONNECTED_1453,SV2V_UNCONNECTED_1454,SV2V_UNCONNECTED_1455,
  SV2V_UNCONNECTED_1456,SV2V_UNCONNECTED_1457,SV2V_UNCONNECTED_1458,
  SV2V_UNCONNECTED_1459,SV2V_UNCONNECTED_1460,SV2V_UNCONNECTED_1461,
  SV2V_UNCONNECTED_1462,SV2V_UNCONNECTED_1463,SV2V_UNCONNECTED_1464,
  SV2V_UNCONNECTED_1465,SV2V_UNCONNECTED_1466,SV2V_UNCONNECTED_1467,SV2V_UNCONNECTED_1468,
  SV2V_UNCONNECTED_1469,SV2V_UNCONNECTED_1470,SV2V_UNCONNECTED_1471,
  SV2V_UNCONNECTED_1472,SV2V_UNCONNECTED_1473,SV2V_UNCONNECTED_1474,
  SV2V_UNCONNECTED_1475,SV2V_UNCONNECTED_1476,SV2V_UNCONNECTED_1477,
  SV2V_UNCONNECTED_1478,SV2V_UNCONNECTED_1479,SV2V_UNCONNECTED_1480,
  SV2V_UNCONNECTED_1481,SV2V_UNCONNECTED_1482,SV2V_UNCONNECTED_1483,
  SV2V_UNCONNECTED_1484,SV2V_UNCONNECTED_1485,SV2V_UNCONNECTED_1486,
  SV2V_UNCONNECTED_1487,SV2V_UNCONNECTED_1488,SV2V_UNCONNECTED_1489,
  SV2V_UNCONNECTED_1490,SV2V_UNCONNECTED_1491,SV2V_UNCONNECTED_1492,
  SV2V_UNCONNECTED_1493,SV2V_UNCONNECTED_1494,SV2V_UNCONNECTED_1495,
  SV2V_UNCONNECTED_1496,SV2V_UNCONNECTED_1497,SV2V_UNCONNECTED_1498,
  SV2V_UNCONNECTED_1499,SV2V_UNCONNECTED_1500,SV2V_UNCONNECTED_1501,
  SV2V_UNCONNECTED_1502,SV2V_UNCONNECTED_1503,SV2V_UNCONNECTED_1504,
  SV2V_UNCONNECTED_1505,SV2V_UNCONNECTED_1506,SV2V_UNCONNECTED_1507,SV2V_UNCONNECTED_1508,
  SV2V_UNCONNECTED_1509,SV2V_UNCONNECTED_1510,SV2V_UNCONNECTED_1511,
  SV2V_UNCONNECTED_1512,SV2V_UNCONNECTED_1513,SV2V_UNCONNECTED_1514,
  SV2V_UNCONNECTED_1515,SV2V_UNCONNECTED_1516,SV2V_UNCONNECTED_1517,
  SV2V_UNCONNECTED_1518,SV2V_UNCONNECTED_1519,SV2V_UNCONNECTED_1520,
  SV2V_UNCONNECTED_1521,SV2V_UNCONNECTED_1522,SV2V_UNCONNECTED_1523,
  SV2V_UNCONNECTED_1524,SV2V_UNCONNECTED_1525,SV2V_UNCONNECTED_1526,
  SV2V_UNCONNECTED_1527,SV2V_UNCONNECTED_1528,SV2V_UNCONNECTED_1529,
  SV2V_UNCONNECTED_1530,SV2V_UNCONNECTED_1531,SV2V_UNCONNECTED_1532,
  SV2V_UNCONNECTED_1533,SV2V_UNCONNECTED_1534,SV2V_UNCONNECTED_1535,
  SV2V_UNCONNECTED_1536,SV2V_UNCONNECTED_1537,SV2V_UNCONNECTED_1538,
  SV2V_UNCONNECTED_1539,SV2V_UNCONNECTED_1540,SV2V_UNCONNECTED_1541,
  SV2V_UNCONNECTED_1542,SV2V_UNCONNECTED_1543,SV2V_UNCONNECTED_1544,
  SV2V_UNCONNECTED_1545,SV2V_UNCONNECTED_1546,SV2V_UNCONNECTED_1547,SV2V_UNCONNECTED_1548,
  SV2V_UNCONNECTED_1549,SV2V_UNCONNECTED_1550,SV2V_UNCONNECTED_1551,
  SV2V_UNCONNECTED_1552,SV2V_UNCONNECTED_1553,SV2V_UNCONNECTED_1554,
  SV2V_UNCONNECTED_1555,SV2V_UNCONNECTED_1556,SV2V_UNCONNECTED_1557,
  SV2V_UNCONNECTED_1558,SV2V_UNCONNECTED_1559,SV2V_UNCONNECTED_1560,
  SV2V_UNCONNECTED_1561,SV2V_UNCONNECTED_1562,SV2V_UNCONNECTED_1563,
  SV2V_UNCONNECTED_1564,SV2V_UNCONNECTED_1565,SV2V_UNCONNECTED_1566,
  SV2V_UNCONNECTED_1567,SV2V_UNCONNECTED_1568,SV2V_UNCONNECTED_1569,
  SV2V_UNCONNECTED_1570,SV2V_UNCONNECTED_1571,SV2V_UNCONNECTED_1572,
  SV2V_UNCONNECTED_1573,SV2V_UNCONNECTED_1574,SV2V_UNCONNECTED_1575,
  SV2V_UNCONNECTED_1576,SV2V_UNCONNECTED_1577,SV2V_UNCONNECTED_1578,
  SV2V_UNCONNECTED_1579,SV2V_UNCONNECTED_1580,SV2V_UNCONNECTED_1581,
  SV2V_UNCONNECTED_1582,SV2V_UNCONNECTED_1583,SV2V_UNCONNECTED_1584,
  SV2V_UNCONNECTED_1585,SV2V_UNCONNECTED_1586,SV2V_UNCONNECTED_1587,SV2V_UNCONNECTED_1588,
  SV2V_UNCONNECTED_1589,SV2V_UNCONNECTED_1590,SV2V_UNCONNECTED_1591,
  SV2V_UNCONNECTED_1592,SV2V_UNCONNECTED_1593,SV2V_UNCONNECTED_1594,
  SV2V_UNCONNECTED_1595,SV2V_UNCONNECTED_1596,SV2V_UNCONNECTED_1597,
  SV2V_UNCONNECTED_1598,SV2V_UNCONNECTED_1599,SV2V_UNCONNECTED_1600,
  SV2V_UNCONNECTED_1601,SV2V_UNCONNECTED_1602,SV2V_UNCONNECTED_1603,
  SV2V_UNCONNECTED_1604,SV2V_UNCONNECTED_1605,SV2V_UNCONNECTED_1606,
  SV2V_UNCONNECTED_1607,SV2V_UNCONNECTED_1608,SV2V_UNCONNECTED_1609,
  SV2V_UNCONNECTED_1610,SV2V_UNCONNECTED_1611,SV2V_UNCONNECTED_1612,
  SV2V_UNCONNECTED_1613,SV2V_UNCONNECTED_1614,SV2V_UNCONNECTED_1615,
  SV2V_UNCONNECTED_1616,SV2V_UNCONNECTED_1617,SV2V_UNCONNECTED_1618,
  SV2V_UNCONNECTED_1619,SV2V_UNCONNECTED_1620,SV2V_UNCONNECTED_1621,
  SV2V_UNCONNECTED_1622,SV2V_UNCONNECTED_1623,SV2V_UNCONNECTED_1624,
  SV2V_UNCONNECTED_1625,SV2V_UNCONNECTED_1626,SV2V_UNCONNECTED_1627,SV2V_UNCONNECTED_1628,
  SV2V_UNCONNECTED_1629,SV2V_UNCONNECTED_1630,SV2V_UNCONNECTED_1631,
  SV2V_UNCONNECTED_1632,SV2V_UNCONNECTED_1633,SV2V_UNCONNECTED_1634,
  SV2V_UNCONNECTED_1635,SV2V_UNCONNECTED_1636,SV2V_UNCONNECTED_1637,
  SV2V_UNCONNECTED_1638,SV2V_UNCONNECTED_1639,SV2V_UNCONNECTED_1640,
  SV2V_UNCONNECTED_1641,SV2V_UNCONNECTED_1642,SV2V_UNCONNECTED_1643,
  SV2V_UNCONNECTED_1644,SV2V_UNCONNECTED_1645,SV2V_UNCONNECTED_1646,
  SV2V_UNCONNECTED_1647,SV2V_UNCONNECTED_1648,SV2V_UNCONNECTED_1649,
  SV2V_UNCONNECTED_1650,SV2V_UNCONNECTED_1651,SV2V_UNCONNECTED_1652,
  SV2V_UNCONNECTED_1653,SV2V_UNCONNECTED_1654,SV2V_UNCONNECTED_1655,
  SV2V_UNCONNECTED_1656,SV2V_UNCONNECTED_1657,SV2V_UNCONNECTED_1658,
  SV2V_UNCONNECTED_1659,SV2V_UNCONNECTED_1660,SV2V_UNCONNECTED_1661,
  SV2V_UNCONNECTED_1662,SV2V_UNCONNECTED_1663,SV2V_UNCONNECTED_1664,
  SV2V_UNCONNECTED_1665,SV2V_UNCONNECTED_1666,SV2V_UNCONNECTED_1667,SV2V_UNCONNECTED_1668,
  SV2V_UNCONNECTED_1669,SV2V_UNCONNECTED_1670,SV2V_UNCONNECTED_1671,
  SV2V_UNCONNECTED_1672,SV2V_UNCONNECTED_1673,SV2V_UNCONNECTED_1674,
  SV2V_UNCONNECTED_1675,SV2V_UNCONNECTED_1676,SV2V_UNCONNECTED_1677,
  SV2V_UNCONNECTED_1678,SV2V_UNCONNECTED_1679,SV2V_UNCONNECTED_1680,
  SV2V_UNCONNECTED_1681,SV2V_UNCONNECTED_1682,SV2V_UNCONNECTED_1683,
  SV2V_UNCONNECTED_1684,SV2V_UNCONNECTED_1685,SV2V_UNCONNECTED_1686,
  SV2V_UNCONNECTED_1687,SV2V_UNCONNECTED_1688,SV2V_UNCONNECTED_1689,
  SV2V_UNCONNECTED_1690,SV2V_UNCONNECTED_1691,SV2V_UNCONNECTED_1692,
  SV2V_UNCONNECTED_1693,SV2V_UNCONNECTED_1694,SV2V_UNCONNECTED_1695,
  SV2V_UNCONNECTED_1696,SV2V_UNCONNECTED_1697,SV2V_UNCONNECTED_1698,
  SV2V_UNCONNECTED_1699,SV2V_UNCONNECTED_1700,SV2V_UNCONNECTED_1701,
  SV2V_UNCONNECTED_1702,SV2V_UNCONNECTED_1703,SV2V_UNCONNECTED_1704,
  SV2V_UNCONNECTED_1705,SV2V_UNCONNECTED_1706,SV2V_UNCONNECTED_1707,SV2V_UNCONNECTED_1708,
  SV2V_UNCONNECTED_1709,SV2V_UNCONNECTED_1710,SV2V_UNCONNECTED_1711,
  SV2V_UNCONNECTED_1712,SV2V_UNCONNECTED_1713,SV2V_UNCONNECTED_1714,
  SV2V_UNCONNECTED_1715,SV2V_UNCONNECTED_1716,SV2V_UNCONNECTED_1717,
  SV2V_UNCONNECTED_1718,SV2V_UNCONNECTED_1719,SV2V_UNCONNECTED_1720,
  SV2V_UNCONNECTED_1721,SV2V_UNCONNECTED_1722,SV2V_UNCONNECTED_1723,
  SV2V_UNCONNECTED_1724,SV2V_UNCONNECTED_1725,SV2V_UNCONNECTED_1726,
  SV2V_UNCONNECTED_1727,SV2V_UNCONNECTED_1728,SV2V_UNCONNECTED_1729,
  SV2V_UNCONNECTED_1730,SV2V_UNCONNECTED_1731,SV2V_UNCONNECTED_1732,
  SV2V_UNCONNECTED_1733,SV2V_UNCONNECTED_1734,SV2V_UNCONNECTED_1735,
  SV2V_UNCONNECTED_1736,SV2V_UNCONNECTED_1737,SV2V_UNCONNECTED_1738,
  SV2V_UNCONNECTED_1739,SV2V_UNCONNECTED_1740,SV2V_UNCONNECTED_1741,
  SV2V_UNCONNECTED_1742,SV2V_UNCONNECTED_1743,SV2V_UNCONNECTED_1744,
  SV2V_UNCONNECTED_1745,SV2V_UNCONNECTED_1746,SV2V_UNCONNECTED_1747,SV2V_UNCONNECTED_1748,
  SV2V_UNCONNECTED_1749,SV2V_UNCONNECTED_1750,SV2V_UNCONNECTED_1751,
  SV2V_UNCONNECTED_1752,SV2V_UNCONNECTED_1753,SV2V_UNCONNECTED_1754,
  SV2V_UNCONNECTED_1755,SV2V_UNCONNECTED_1756,SV2V_UNCONNECTED_1757,
  SV2V_UNCONNECTED_1758,SV2V_UNCONNECTED_1759,SV2V_UNCONNECTED_1760,
  SV2V_UNCONNECTED_1761,SV2V_UNCONNECTED_1762,SV2V_UNCONNECTED_1763,
  SV2V_UNCONNECTED_1764,SV2V_UNCONNECTED_1765,SV2V_UNCONNECTED_1766,
  SV2V_UNCONNECTED_1767,SV2V_UNCONNECTED_1768,SV2V_UNCONNECTED_1769,
  SV2V_UNCONNECTED_1770,SV2V_UNCONNECTED_1771,SV2V_UNCONNECTED_1772,
  SV2V_UNCONNECTED_1773,SV2V_UNCONNECTED_1774,SV2V_UNCONNECTED_1775,
  SV2V_UNCONNECTED_1776,SV2V_UNCONNECTED_1777,SV2V_UNCONNECTED_1778,
  SV2V_UNCONNECTED_1779,SV2V_UNCONNECTED_1780,SV2V_UNCONNECTED_1781,
  SV2V_UNCONNECTED_1782,SV2V_UNCONNECTED_1783,SV2V_UNCONNECTED_1784,
  SV2V_UNCONNECTED_1785,SV2V_UNCONNECTED_1786,SV2V_UNCONNECTED_1787,SV2V_UNCONNECTED_1788,
  SV2V_UNCONNECTED_1789,SV2V_UNCONNECTED_1790,SV2V_UNCONNECTED_1791,
  SV2V_UNCONNECTED_1792,SV2V_UNCONNECTED_1793,SV2V_UNCONNECTED_1794,
  SV2V_UNCONNECTED_1795,SV2V_UNCONNECTED_1796,SV2V_UNCONNECTED_1797,
  SV2V_UNCONNECTED_1798,SV2V_UNCONNECTED_1799,SV2V_UNCONNECTED_1800,
  SV2V_UNCONNECTED_1801,SV2V_UNCONNECTED_1802,SV2V_UNCONNECTED_1803,
  SV2V_UNCONNECTED_1804,SV2V_UNCONNECTED_1805,SV2V_UNCONNECTED_1806,
  SV2V_UNCONNECTED_1807,SV2V_UNCONNECTED_1808,SV2V_UNCONNECTED_1809,
  SV2V_UNCONNECTED_1810,SV2V_UNCONNECTED_1811,SV2V_UNCONNECTED_1812,
  SV2V_UNCONNECTED_1813,SV2V_UNCONNECTED_1814,SV2V_UNCONNECTED_1815,
  SV2V_UNCONNECTED_1816,SV2V_UNCONNECTED_1817,SV2V_UNCONNECTED_1818,
  SV2V_UNCONNECTED_1819,SV2V_UNCONNECTED_1820,SV2V_UNCONNECTED_1821,
  SV2V_UNCONNECTED_1822,SV2V_UNCONNECTED_1823,SV2V_UNCONNECTED_1824,
  SV2V_UNCONNECTED_1825,SV2V_UNCONNECTED_1826,SV2V_UNCONNECTED_1827,SV2V_UNCONNECTED_1828,
  SV2V_UNCONNECTED_1829,SV2V_UNCONNECTED_1830,SV2V_UNCONNECTED_1831,
  SV2V_UNCONNECTED_1832,SV2V_UNCONNECTED_1833,SV2V_UNCONNECTED_1834,
  SV2V_UNCONNECTED_1835,SV2V_UNCONNECTED_1836,SV2V_UNCONNECTED_1837,
  SV2V_UNCONNECTED_1838,SV2V_UNCONNECTED_1839,SV2V_UNCONNECTED_1840,
  SV2V_UNCONNECTED_1841,SV2V_UNCONNECTED_1842,SV2V_UNCONNECTED_1843,
  SV2V_UNCONNECTED_1844,SV2V_UNCONNECTED_1845,SV2V_UNCONNECTED_1846,
  SV2V_UNCONNECTED_1847,SV2V_UNCONNECTED_1848,SV2V_UNCONNECTED_1849,
  SV2V_UNCONNECTED_1850,SV2V_UNCONNECTED_1851,SV2V_UNCONNECTED_1852,
  SV2V_UNCONNECTED_1853,SV2V_UNCONNECTED_1854,SV2V_UNCONNECTED_1855,
  SV2V_UNCONNECTED_1856,SV2V_UNCONNECTED_1857,SV2V_UNCONNECTED_1858,
  SV2V_UNCONNECTED_1859,SV2V_UNCONNECTED_1860,SV2V_UNCONNECTED_1861,
  SV2V_UNCONNECTED_1862,SV2V_UNCONNECTED_1863,SV2V_UNCONNECTED_1864,
  SV2V_UNCONNECTED_1865,SV2V_UNCONNECTED_1866,SV2V_UNCONNECTED_1867,SV2V_UNCONNECTED_1868,
  SV2V_UNCONNECTED_1869,SV2V_UNCONNECTED_1870,SV2V_UNCONNECTED_1871,
  SV2V_UNCONNECTED_1872,SV2V_UNCONNECTED_1873,SV2V_UNCONNECTED_1874,
  SV2V_UNCONNECTED_1875,SV2V_UNCONNECTED_1876,SV2V_UNCONNECTED_1877,
  SV2V_UNCONNECTED_1878,SV2V_UNCONNECTED_1879,SV2V_UNCONNECTED_1880,
  SV2V_UNCONNECTED_1881,SV2V_UNCONNECTED_1882,SV2V_UNCONNECTED_1883,
  SV2V_UNCONNECTED_1884,SV2V_UNCONNECTED_1885,SV2V_UNCONNECTED_1886,
  SV2V_UNCONNECTED_1887,SV2V_UNCONNECTED_1888,SV2V_UNCONNECTED_1889,
  SV2V_UNCONNECTED_1890,SV2V_UNCONNECTED_1891,SV2V_UNCONNECTED_1892,
  SV2V_UNCONNECTED_1893,SV2V_UNCONNECTED_1894,SV2V_UNCONNECTED_1895,
  SV2V_UNCONNECTED_1896,SV2V_UNCONNECTED_1897,SV2V_UNCONNECTED_1898,
  SV2V_UNCONNECTED_1899,SV2V_UNCONNECTED_1900,SV2V_UNCONNECTED_1901,
  SV2V_UNCONNECTED_1902,SV2V_UNCONNECTED_1903,SV2V_UNCONNECTED_1904,
  SV2V_UNCONNECTED_1905,SV2V_UNCONNECTED_1906,SV2V_UNCONNECTED_1907,SV2V_UNCONNECTED_1908,
  SV2V_UNCONNECTED_1909,SV2V_UNCONNECTED_1910,SV2V_UNCONNECTED_1911,
  SV2V_UNCONNECTED_1912,SV2V_UNCONNECTED_1913,SV2V_UNCONNECTED_1914,
  SV2V_UNCONNECTED_1915,SV2V_UNCONNECTED_1916,SV2V_UNCONNECTED_1917,
  SV2V_UNCONNECTED_1918,SV2V_UNCONNECTED_1919,SV2V_UNCONNECTED_1920,
  SV2V_UNCONNECTED_1921,SV2V_UNCONNECTED_1922,SV2V_UNCONNECTED_1923,
  SV2V_UNCONNECTED_1924,SV2V_UNCONNECTED_1925,SV2V_UNCONNECTED_1926,
  SV2V_UNCONNECTED_1927,SV2V_UNCONNECTED_1928,SV2V_UNCONNECTED_1929,
  SV2V_UNCONNECTED_1930,SV2V_UNCONNECTED_1931,SV2V_UNCONNECTED_1932,
  SV2V_UNCONNECTED_1933,SV2V_UNCONNECTED_1934,SV2V_UNCONNECTED_1935,
  SV2V_UNCONNECTED_1936,SV2V_UNCONNECTED_1937,SV2V_UNCONNECTED_1938,
  SV2V_UNCONNECTED_1939,SV2V_UNCONNECTED_1940,SV2V_UNCONNECTED_1941,
  SV2V_UNCONNECTED_1942,SV2V_UNCONNECTED_1943,SV2V_UNCONNECTED_1944,
  SV2V_UNCONNECTED_1945,SV2V_UNCONNECTED_1946,SV2V_UNCONNECTED_1947,SV2V_UNCONNECTED_1948,
  SV2V_UNCONNECTED_1949,SV2V_UNCONNECTED_1950,SV2V_UNCONNECTED_1951,
  SV2V_UNCONNECTED_1952,SV2V_UNCONNECTED_1953,SV2V_UNCONNECTED_1954,
  SV2V_UNCONNECTED_1955,SV2V_UNCONNECTED_1956,SV2V_UNCONNECTED_1957,
  SV2V_UNCONNECTED_1958,SV2V_UNCONNECTED_1959,SV2V_UNCONNECTED_1960,
  SV2V_UNCONNECTED_1961,SV2V_UNCONNECTED_1962,SV2V_UNCONNECTED_1963,
  SV2V_UNCONNECTED_1964,SV2V_UNCONNECTED_1965,SV2V_UNCONNECTED_1966,
  SV2V_UNCONNECTED_1967,SV2V_UNCONNECTED_1968,SV2V_UNCONNECTED_1969,
  SV2V_UNCONNECTED_1970,SV2V_UNCONNECTED_1971,SV2V_UNCONNECTED_1972,
  SV2V_UNCONNECTED_1973,SV2V_UNCONNECTED_1974,SV2V_UNCONNECTED_1975,
  SV2V_UNCONNECTED_1976,SV2V_UNCONNECTED_1977,SV2V_UNCONNECTED_1978,
  SV2V_UNCONNECTED_1979,SV2V_UNCONNECTED_1980,SV2V_UNCONNECTED_1981,
  SV2V_UNCONNECTED_1982,SV2V_UNCONNECTED_1983,SV2V_UNCONNECTED_1984,
  SV2V_UNCONNECTED_1985,SV2V_UNCONNECTED_1986,SV2V_UNCONNECTED_1987,SV2V_UNCONNECTED_1988,
  SV2V_UNCONNECTED_1989,SV2V_UNCONNECTED_1990,SV2V_UNCONNECTED_1991,
  SV2V_UNCONNECTED_1992,SV2V_UNCONNECTED_1993,SV2V_UNCONNECTED_1994,
  SV2V_UNCONNECTED_1995,SV2V_UNCONNECTED_1996,SV2V_UNCONNECTED_1997,
  SV2V_UNCONNECTED_1998,SV2V_UNCONNECTED_1999,SV2V_UNCONNECTED_2000,
  SV2V_UNCONNECTED_2001,SV2V_UNCONNECTED_2002,SV2V_UNCONNECTED_2003,
  SV2V_UNCONNECTED_2004,SV2V_UNCONNECTED_2005,SV2V_UNCONNECTED_2006,
  SV2V_UNCONNECTED_2007,SV2V_UNCONNECTED_2008,SV2V_UNCONNECTED_2009,
  SV2V_UNCONNECTED_2010,SV2V_UNCONNECTED_2011,SV2V_UNCONNECTED_2012,
  SV2V_UNCONNECTED_2013,SV2V_UNCONNECTED_2014,SV2V_UNCONNECTED_2015,
  SV2V_UNCONNECTED_2016,SV2V_UNCONNECTED_2017,SV2V_UNCONNECTED_2018,
  SV2V_UNCONNECTED_2019,SV2V_UNCONNECTED_2020,SV2V_UNCONNECTED_2021,
  SV2V_UNCONNECTED_2022,SV2V_UNCONNECTED_2023,SV2V_UNCONNECTED_2024,
  SV2V_UNCONNECTED_2025,SV2V_UNCONNECTED_2026,SV2V_UNCONNECTED_2027,SV2V_UNCONNECTED_2028,
  SV2V_UNCONNECTED_2029,SV2V_UNCONNECTED_2030,SV2V_UNCONNECTED_2031,
  SV2V_UNCONNECTED_2032,SV2V_UNCONNECTED_2033,SV2V_UNCONNECTED_2034,
  SV2V_UNCONNECTED_2035,SV2V_UNCONNECTED_2036,SV2V_UNCONNECTED_2037,
  SV2V_UNCONNECTED_2038,SV2V_UNCONNECTED_2039,SV2V_UNCONNECTED_2040,
  SV2V_UNCONNECTED_2041,SV2V_UNCONNECTED_2042,SV2V_UNCONNECTED_2043,
  SV2V_UNCONNECTED_2044,SV2V_UNCONNECTED_2045,SV2V_UNCONNECTED_2046,
  SV2V_UNCONNECTED_2047,SV2V_UNCONNECTED_2048,SV2V_UNCONNECTED_2049,
  SV2V_UNCONNECTED_2050,SV2V_UNCONNECTED_2051,SV2V_UNCONNECTED_2052,
  SV2V_UNCONNECTED_2053,SV2V_UNCONNECTED_2054,SV2V_UNCONNECTED_2055,
  SV2V_UNCONNECTED_2056,SV2V_UNCONNECTED_2057,SV2V_UNCONNECTED_2058,
  SV2V_UNCONNECTED_2059,SV2V_UNCONNECTED_2060,SV2V_UNCONNECTED_2061,
  SV2V_UNCONNECTED_2062,SV2V_UNCONNECTED_2063,SV2V_UNCONNECTED_2064,
  SV2V_UNCONNECTED_2065,SV2V_UNCONNECTED_2066,SV2V_UNCONNECTED_2067,SV2V_UNCONNECTED_2068,
  SV2V_UNCONNECTED_2069,SV2V_UNCONNECTED_2070,SV2V_UNCONNECTED_2071,
  SV2V_UNCONNECTED_2072,SV2V_UNCONNECTED_2073,SV2V_UNCONNECTED_2074,
  SV2V_UNCONNECTED_2075,SV2V_UNCONNECTED_2076,SV2V_UNCONNECTED_2077,
  SV2V_UNCONNECTED_2078,SV2V_UNCONNECTED_2079,SV2V_UNCONNECTED_2080,
  SV2V_UNCONNECTED_2081,SV2V_UNCONNECTED_2082,SV2V_UNCONNECTED_2083,
  SV2V_UNCONNECTED_2084,SV2V_UNCONNECTED_2085,SV2V_UNCONNECTED_2086,
  SV2V_UNCONNECTED_2087,SV2V_UNCONNECTED_2088,SV2V_UNCONNECTED_2089,
  SV2V_UNCONNECTED_2090,SV2V_UNCONNECTED_2091,SV2V_UNCONNECTED_2092,
  SV2V_UNCONNECTED_2093,SV2V_UNCONNECTED_2094,SV2V_UNCONNECTED_2095,
  SV2V_UNCONNECTED_2096,SV2V_UNCONNECTED_2097,SV2V_UNCONNECTED_2098,
  SV2V_UNCONNECTED_2099,SV2V_UNCONNECTED_2100,SV2V_UNCONNECTED_2101,
  SV2V_UNCONNECTED_2102,SV2V_UNCONNECTED_2103,SV2V_UNCONNECTED_2104,
  SV2V_UNCONNECTED_2105,SV2V_UNCONNECTED_2106,SV2V_UNCONNECTED_2107,SV2V_UNCONNECTED_2108,
  SV2V_UNCONNECTED_2109,SV2V_UNCONNECTED_2110,SV2V_UNCONNECTED_2111,
  SV2V_UNCONNECTED_2112,SV2V_UNCONNECTED_2113,SV2V_UNCONNECTED_2114,
  SV2V_UNCONNECTED_2115,SV2V_UNCONNECTED_2116,SV2V_UNCONNECTED_2117,
  SV2V_UNCONNECTED_2118,SV2V_UNCONNECTED_2119,SV2V_UNCONNECTED_2120,
  SV2V_UNCONNECTED_2121,SV2V_UNCONNECTED_2122,SV2V_UNCONNECTED_2123,
  SV2V_UNCONNECTED_2124,SV2V_UNCONNECTED_2125,SV2V_UNCONNECTED_2126,
  SV2V_UNCONNECTED_2127,SV2V_UNCONNECTED_2128,SV2V_UNCONNECTED_2129,
  SV2V_UNCONNECTED_2130,SV2V_UNCONNECTED_2131,SV2V_UNCONNECTED_2132,
  SV2V_UNCONNECTED_2133,SV2V_UNCONNECTED_2134,SV2V_UNCONNECTED_2135,
  SV2V_UNCONNECTED_2136,SV2V_UNCONNECTED_2137,SV2V_UNCONNECTED_2138,
  SV2V_UNCONNECTED_2139,SV2V_UNCONNECTED_2140,SV2V_UNCONNECTED_2141,
  SV2V_UNCONNECTED_2142,SV2V_UNCONNECTED_2143,SV2V_UNCONNECTED_2144,
  SV2V_UNCONNECTED_2145,SV2V_UNCONNECTED_2146,SV2V_UNCONNECTED_2147,SV2V_UNCONNECTED_2148,
  SV2V_UNCONNECTED_2149,SV2V_UNCONNECTED_2150,SV2V_UNCONNECTED_2151,
  SV2V_UNCONNECTED_2152,SV2V_UNCONNECTED_2153,SV2V_UNCONNECTED_2154,
  SV2V_UNCONNECTED_2155,SV2V_UNCONNECTED_2156,SV2V_UNCONNECTED_2157,
  SV2V_UNCONNECTED_2158,SV2V_UNCONNECTED_2159,SV2V_UNCONNECTED_2160,
  SV2V_UNCONNECTED_2161,SV2V_UNCONNECTED_2162,SV2V_UNCONNECTED_2163,
  SV2V_UNCONNECTED_2164,SV2V_UNCONNECTED_2165,SV2V_UNCONNECTED_2166,
  SV2V_UNCONNECTED_2167,SV2V_UNCONNECTED_2168,SV2V_UNCONNECTED_2169,
  SV2V_UNCONNECTED_2170,SV2V_UNCONNECTED_2171,SV2V_UNCONNECTED_2172,
  SV2V_UNCONNECTED_2173,SV2V_UNCONNECTED_2174,SV2V_UNCONNECTED_2175,
  SV2V_UNCONNECTED_2176,SV2V_UNCONNECTED_2177,SV2V_UNCONNECTED_2178,
  SV2V_UNCONNECTED_2179,SV2V_UNCONNECTED_2180,SV2V_UNCONNECTED_2181,
  SV2V_UNCONNECTED_2182,SV2V_UNCONNECTED_2183,SV2V_UNCONNECTED_2184,
  SV2V_UNCONNECTED_2185,SV2V_UNCONNECTED_2186,SV2V_UNCONNECTED_2187,SV2V_UNCONNECTED_2188,
  SV2V_UNCONNECTED_2189,SV2V_UNCONNECTED_2190,SV2V_UNCONNECTED_2191,
  SV2V_UNCONNECTED_2192,SV2V_UNCONNECTED_2193,SV2V_UNCONNECTED_2194,
  SV2V_UNCONNECTED_2195,SV2V_UNCONNECTED_2196,SV2V_UNCONNECTED_2197,
  SV2V_UNCONNECTED_2198,SV2V_UNCONNECTED_2199,SV2V_UNCONNECTED_2200,
  SV2V_UNCONNECTED_2201,SV2V_UNCONNECTED_2202,SV2V_UNCONNECTED_2203,
  SV2V_UNCONNECTED_2204,SV2V_UNCONNECTED_2205,SV2V_UNCONNECTED_2206,
  SV2V_UNCONNECTED_2207,SV2V_UNCONNECTED_2208,SV2V_UNCONNECTED_2209,
  SV2V_UNCONNECTED_2210,SV2V_UNCONNECTED_2211,SV2V_UNCONNECTED_2212,
  SV2V_UNCONNECTED_2213,SV2V_UNCONNECTED_2214,SV2V_UNCONNECTED_2215,
  SV2V_UNCONNECTED_2216,SV2V_UNCONNECTED_2217,SV2V_UNCONNECTED_2218,
  SV2V_UNCONNECTED_2219,SV2V_UNCONNECTED_2220,SV2V_UNCONNECTED_2221,
  SV2V_UNCONNECTED_2222,SV2V_UNCONNECTED_2223,SV2V_UNCONNECTED_2224,
  SV2V_UNCONNECTED_2225,SV2V_UNCONNECTED_2226,SV2V_UNCONNECTED_2227,SV2V_UNCONNECTED_2228,
  SV2V_UNCONNECTED_2229,SV2V_UNCONNECTED_2230,SV2V_UNCONNECTED_2231,
  SV2V_UNCONNECTED_2232,SV2V_UNCONNECTED_2233,SV2V_UNCONNECTED_2234,
  SV2V_UNCONNECTED_2235,SV2V_UNCONNECTED_2236,SV2V_UNCONNECTED_2237,
  SV2V_UNCONNECTED_2238,SV2V_UNCONNECTED_2239,SV2V_UNCONNECTED_2240,
  SV2V_UNCONNECTED_2241,SV2V_UNCONNECTED_2242,SV2V_UNCONNECTED_2243,
  SV2V_UNCONNECTED_2244,SV2V_UNCONNECTED_2245,SV2V_UNCONNECTED_2246,
  SV2V_UNCONNECTED_2247,SV2V_UNCONNECTED_2248,SV2V_UNCONNECTED_2249,
  SV2V_UNCONNECTED_2250,SV2V_UNCONNECTED_2251,SV2V_UNCONNECTED_2252,
  SV2V_UNCONNECTED_2253,SV2V_UNCONNECTED_2254,SV2V_UNCONNECTED_2255,
  SV2V_UNCONNECTED_2256,SV2V_UNCONNECTED_2257,SV2V_UNCONNECTED_2258,
  SV2V_UNCONNECTED_2259,SV2V_UNCONNECTED_2260,SV2V_UNCONNECTED_2261,
  SV2V_UNCONNECTED_2262,SV2V_UNCONNECTED_2263,SV2V_UNCONNECTED_2264,
  SV2V_UNCONNECTED_2265,SV2V_UNCONNECTED_2266,SV2V_UNCONNECTED_2267,SV2V_UNCONNECTED_2268,
  SV2V_UNCONNECTED_2269,SV2V_UNCONNECTED_2270,SV2V_UNCONNECTED_2271,
  SV2V_UNCONNECTED_2272,SV2V_UNCONNECTED_2273,SV2V_UNCONNECTED_2274,
  SV2V_UNCONNECTED_2275,SV2V_UNCONNECTED_2276,SV2V_UNCONNECTED_2277,
  SV2V_UNCONNECTED_2278,SV2V_UNCONNECTED_2279,SV2V_UNCONNECTED_2280,
  SV2V_UNCONNECTED_2281,SV2V_UNCONNECTED_2282,SV2V_UNCONNECTED_2283,
  SV2V_UNCONNECTED_2284,SV2V_UNCONNECTED_2285,SV2V_UNCONNECTED_2286,
  SV2V_UNCONNECTED_2287,SV2V_UNCONNECTED_2288,SV2V_UNCONNECTED_2289,
  SV2V_UNCONNECTED_2290,SV2V_UNCONNECTED_2291,SV2V_UNCONNECTED_2292,
  SV2V_UNCONNECTED_2293,SV2V_UNCONNECTED_2294,SV2V_UNCONNECTED_2295,
  SV2V_UNCONNECTED_2296,SV2V_UNCONNECTED_2297,SV2V_UNCONNECTED_2298,
  SV2V_UNCONNECTED_2299,SV2V_UNCONNECTED_2300,SV2V_UNCONNECTED_2301,
  SV2V_UNCONNECTED_2302,SV2V_UNCONNECTED_2303,SV2V_UNCONNECTED_2304,
  SV2V_UNCONNECTED_2305,SV2V_UNCONNECTED_2306,SV2V_UNCONNECTED_2307,SV2V_UNCONNECTED_2308,
  SV2V_UNCONNECTED_2309,SV2V_UNCONNECTED_2310,SV2V_UNCONNECTED_2311,
  SV2V_UNCONNECTED_2312,SV2V_UNCONNECTED_2313,SV2V_UNCONNECTED_2314,
  SV2V_UNCONNECTED_2315,SV2V_UNCONNECTED_2316,SV2V_UNCONNECTED_2317,
  SV2V_UNCONNECTED_2318,SV2V_UNCONNECTED_2319,SV2V_UNCONNECTED_2320,
  SV2V_UNCONNECTED_2321,SV2V_UNCONNECTED_2322,SV2V_UNCONNECTED_2323,
  SV2V_UNCONNECTED_2324,SV2V_UNCONNECTED_2325,SV2V_UNCONNECTED_2326,
  SV2V_UNCONNECTED_2327,SV2V_UNCONNECTED_2328,SV2V_UNCONNECTED_2329,
  SV2V_UNCONNECTED_2330,SV2V_UNCONNECTED_2331,SV2V_UNCONNECTED_2332,
  SV2V_UNCONNECTED_2333,SV2V_UNCONNECTED_2334,SV2V_UNCONNECTED_2335,
  SV2V_UNCONNECTED_2336,SV2V_UNCONNECTED_2337,SV2V_UNCONNECTED_2338,
  SV2V_UNCONNECTED_2339,SV2V_UNCONNECTED_2340,SV2V_UNCONNECTED_2341,
  SV2V_UNCONNECTED_2342,SV2V_UNCONNECTED_2343,SV2V_UNCONNECTED_2344,
  SV2V_UNCONNECTED_2345,SV2V_UNCONNECTED_2346,SV2V_UNCONNECTED_2347,SV2V_UNCONNECTED_2348,
  SV2V_UNCONNECTED_2349,SV2V_UNCONNECTED_2350,SV2V_UNCONNECTED_2351,
  SV2V_UNCONNECTED_2352,SV2V_UNCONNECTED_2353,SV2V_UNCONNECTED_2354,
  SV2V_UNCONNECTED_2355,SV2V_UNCONNECTED_2356,SV2V_UNCONNECTED_2357,
  SV2V_UNCONNECTED_2358,SV2V_UNCONNECTED_2359,SV2V_UNCONNECTED_2360,
  SV2V_UNCONNECTED_2361,SV2V_UNCONNECTED_2362,SV2V_UNCONNECTED_2363,
  SV2V_UNCONNECTED_2364,SV2V_UNCONNECTED_2365,SV2V_UNCONNECTED_2366,
  SV2V_UNCONNECTED_2367,SV2V_UNCONNECTED_2368,SV2V_UNCONNECTED_2369,
  SV2V_UNCONNECTED_2370,SV2V_UNCONNECTED_2371,SV2V_UNCONNECTED_2372,
  SV2V_UNCONNECTED_2373,SV2V_UNCONNECTED_2374,SV2V_UNCONNECTED_2375,
  SV2V_UNCONNECTED_2376,SV2V_UNCONNECTED_2377,SV2V_UNCONNECTED_2378,
  SV2V_UNCONNECTED_2379,SV2V_UNCONNECTED_2380,SV2V_UNCONNECTED_2381,
  SV2V_UNCONNECTED_2382,SV2V_UNCONNECTED_2383,SV2V_UNCONNECTED_2384,
  SV2V_UNCONNECTED_2385,SV2V_UNCONNECTED_2386,SV2V_UNCONNECTED_2387,SV2V_UNCONNECTED_2388,
  SV2V_UNCONNECTED_2389,SV2V_UNCONNECTED_2390,SV2V_UNCONNECTED_2391,
  SV2V_UNCONNECTED_2392,SV2V_UNCONNECTED_2393,SV2V_UNCONNECTED_2394,
  SV2V_UNCONNECTED_2395,SV2V_UNCONNECTED_2396,SV2V_UNCONNECTED_2397,
  SV2V_UNCONNECTED_2398,SV2V_UNCONNECTED_2399,SV2V_UNCONNECTED_2400,
  SV2V_UNCONNECTED_2401,SV2V_UNCONNECTED_2402,SV2V_UNCONNECTED_2403,
  SV2V_UNCONNECTED_2404,SV2V_UNCONNECTED_2405,SV2V_UNCONNECTED_2406,
  SV2V_UNCONNECTED_2407,SV2V_UNCONNECTED_2408,SV2V_UNCONNECTED_2409,
  SV2V_UNCONNECTED_2410,SV2V_UNCONNECTED_2411,SV2V_UNCONNECTED_2412,
  SV2V_UNCONNECTED_2413,SV2V_UNCONNECTED_2414,SV2V_UNCONNECTED_2415,
  SV2V_UNCONNECTED_2416,SV2V_UNCONNECTED_2417,SV2V_UNCONNECTED_2418,
  SV2V_UNCONNECTED_2419,SV2V_UNCONNECTED_2420,SV2V_UNCONNECTED_2421,
  SV2V_UNCONNECTED_2422,SV2V_UNCONNECTED_2423,SV2V_UNCONNECTED_2424,
  SV2V_UNCONNECTED_2425,SV2V_UNCONNECTED_2426,SV2V_UNCONNECTED_2427,SV2V_UNCONNECTED_2428,
  SV2V_UNCONNECTED_2429,SV2V_UNCONNECTED_2430,SV2V_UNCONNECTED_2431,
  SV2V_UNCONNECTED_2432,SV2V_UNCONNECTED_2433,SV2V_UNCONNECTED_2434,
  SV2V_UNCONNECTED_2435,SV2V_UNCONNECTED_2436,SV2V_UNCONNECTED_2437,
  SV2V_UNCONNECTED_2438,SV2V_UNCONNECTED_2439,SV2V_UNCONNECTED_2440,
  SV2V_UNCONNECTED_2441,SV2V_UNCONNECTED_2442,SV2V_UNCONNECTED_2443,
  SV2V_UNCONNECTED_2444,SV2V_UNCONNECTED_2445,SV2V_UNCONNECTED_2446,
  SV2V_UNCONNECTED_2447,SV2V_UNCONNECTED_2448,SV2V_UNCONNECTED_2449,
  SV2V_UNCONNECTED_2450,SV2V_UNCONNECTED_2451,SV2V_UNCONNECTED_2452,
  SV2V_UNCONNECTED_2453,SV2V_UNCONNECTED_2454,SV2V_UNCONNECTED_2455,
  SV2V_UNCONNECTED_2456,SV2V_UNCONNECTED_2457,SV2V_UNCONNECTED_2458,
  SV2V_UNCONNECTED_2459,SV2V_UNCONNECTED_2460,SV2V_UNCONNECTED_2461,
  SV2V_UNCONNECTED_2462,SV2V_UNCONNECTED_2463,SV2V_UNCONNECTED_2464,
  SV2V_UNCONNECTED_2465,SV2V_UNCONNECTED_2466,SV2V_UNCONNECTED_2467,SV2V_UNCONNECTED_2468,
  SV2V_UNCONNECTED_2469,SV2V_UNCONNECTED_2470,SV2V_UNCONNECTED_2471,
  SV2V_UNCONNECTED_2472,SV2V_UNCONNECTED_2473,SV2V_UNCONNECTED_2474,
  SV2V_UNCONNECTED_2475,SV2V_UNCONNECTED_2476,SV2V_UNCONNECTED_2477,
  SV2V_UNCONNECTED_2478,SV2V_UNCONNECTED_2479,SV2V_UNCONNECTED_2480,
  SV2V_UNCONNECTED_2481,SV2V_UNCONNECTED_2482,SV2V_UNCONNECTED_2483,
  SV2V_UNCONNECTED_2484,SV2V_UNCONNECTED_2485,SV2V_UNCONNECTED_2486,
  SV2V_UNCONNECTED_2487,SV2V_UNCONNECTED_2488,SV2V_UNCONNECTED_2489,
  SV2V_UNCONNECTED_2490,SV2V_UNCONNECTED_2491,SV2V_UNCONNECTED_2492,
  SV2V_UNCONNECTED_2493,SV2V_UNCONNECTED_2494,SV2V_UNCONNECTED_2495,
  SV2V_UNCONNECTED_2496,SV2V_UNCONNECTED_2497,SV2V_UNCONNECTED_2498,
  SV2V_UNCONNECTED_2499,SV2V_UNCONNECTED_2500,SV2V_UNCONNECTED_2501,
  SV2V_UNCONNECTED_2502,SV2V_UNCONNECTED_2503,SV2V_UNCONNECTED_2504,
  SV2V_UNCONNECTED_2505,SV2V_UNCONNECTED_2506,SV2V_UNCONNECTED_2507,SV2V_UNCONNECTED_2508,
  SV2V_UNCONNECTED_2509,SV2V_UNCONNECTED_2510,SV2V_UNCONNECTED_2511,
  SV2V_UNCONNECTED_2512,SV2V_UNCONNECTED_2513,SV2V_UNCONNECTED_2514,
  SV2V_UNCONNECTED_2515,SV2V_UNCONNECTED_2516,SV2V_UNCONNECTED_2517,
  SV2V_UNCONNECTED_2518,SV2V_UNCONNECTED_2519,SV2V_UNCONNECTED_2520,
  SV2V_UNCONNECTED_2521,SV2V_UNCONNECTED_2522,SV2V_UNCONNECTED_2523,
  SV2V_UNCONNECTED_2524,SV2V_UNCONNECTED_2525,SV2V_UNCONNECTED_2526,
  SV2V_UNCONNECTED_2527,SV2V_UNCONNECTED_2528,SV2V_UNCONNECTED_2529,
  SV2V_UNCONNECTED_2530,SV2V_UNCONNECTED_2531,SV2V_UNCONNECTED_2532,
  SV2V_UNCONNECTED_2533,SV2V_UNCONNECTED_2534,SV2V_UNCONNECTED_2535,
  SV2V_UNCONNECTED_2536,SV2V_UNCONNECTED_2537,SV2V_UNCONNECTED_2538,
  SV2V_UNCONNECTED_2539,SV2V_UNCONNECTED_2540,SV2V_UNCONNECTED_2541,
  SV2V_UNCONNECTED_2542,SV2V_UNCONNECTED_2543,SV2V_UNCONNECTED_2544,
  SV2V_UNCONNECTED_2545,SV2V_UNCONNECTED_2546,SV2V_UNCONNECTED_2547,SV2V_UNCONNECTED_2548,
  SV2V_UNCONNECTED_2549,SV2V_UNCONNECTED_2550,SV2V_UNCONNECTED_2551,
  SV2V_UNCONNECTED_2552,SV2V_UNCONNECTED_2553,SV2V_UNCONNECTED_2554,
  SV2V_UNCONNECTED_2555,SV2V_UNCONNECTED_2556,SV2V_UNCONNECTED_2557,
  SV2V_UNCONNECTED_2558,SV2V_UNCONNECTED_2559,SV2V_UNCONNECTED_2560,
  SV2V_UNCONNECTED_2561,SV2V_UNCONNECTED_2562,SV2V_UNCONNECTED_2563,
  SV2V_UNCONNECTED_2564,SV2V_UNCONNECTED_2565,SV2V_UNCONNECTED_2566,
  SV2V_UNCONNECTED_2567,SV2V_UNCONNECTED_2568,SV2V_UNCONNECTED_2569,
  SV2V_UNCONNECTED_2570,SV2V_UNCONNECTED_2571,SV2V_UNCONNECTED_2572,
  SV2V_UNCONNECTED_2573,SV2V_UNCONNECTED_2574,SV2V_UNCONNECTED_2575,
  SV2V_UNCONNECTED_2576,SV2V_UNCONNECTED_2577,SV2V_UNCONNECTED_2578,
  SV2V_UNCONNECTED_2579,SV2V_UNCONNECTED_2580,SV2V_UNCONNECTED_2581,
  SV2V_UNCONNECTED_2582,SV2V_UNCONNECTED_2583,SV2V_UNCONNECTED_2584,
  SV2V_UNCONNECTED_2585,SV2V_UNCONNECTED_2586,SV2V_UNCONNECTED_2587,SV2V_UNCONNECTED_2588,
  SV2V_UNCONNECTED_2589,SV2V_UNCONNECTED_2590,SV2V_UNCONNECTED_2591,
  SV2V_UNCONNECTED_2592,SV2V_UNCONNECTED_2593,SV2V_UNCONNECTED_2594,
  SV2V_UNCONNECTED_2595,SV2V_UNCONNECTED_2596,SV2V_UNCONNECTED_2597,
  SV2V_UNCONNECTED_2598,SV2V_UNCONNECTED_2599,SV2V_UNCONNECTED_2600,
  SV2V_UNCONNECTED_2601,SV2V_UNCONNECTED_2602,SV2V_UNCONNECTED_2603,
  SV2V_UNCONNECTED_2604,SV2V_UNCONNECTED_2605,SV2V_UNCONNECTED_2606,
  SV2V_UNCONNECTED_2607,SV2V_UNCONNECTED_2608,SV2V_UNCONNECTED_2609,
  SV2V_UNCONNECTED_2610,SV2V_UNCONNECTED_2611,SV2V_UNCONNECTED_2612,
  SV2V_UNCONNECTED_2613,SV2V_UNCONNECTED_2614,SV2V_UNCONNECTED_2615,
  SV2V_UNCONNECTED_2616,SV2V_UNCONNECTED_2617,SV2V_UNCONNECTED_2618,
  SV2V_UNCONNECTED_2619,SV2V_UNCONNECTED_2620,SV2V_UNCONNECTED_2621,
  SV2V_UNCONNECTED_2622,SV2V_UNCONNECTED_2623,SV2V_UNCONNECTED_2624,
  SV2V_UNCONNECTED_2625,SV2V_UNCONNECTED_2626,SV2V_UNCONNECTED_2627,SV2V_UNCONNECTED_2628,
  SV2V_UNCONNECTED_2629,SV2V_UNCONNECTED_2630,SV2V_UNCONNECTED_2631,
  SV2V_UNCONNECTED_2632,SV2V_UNCONNECTED_2633,SV2V_UNCONNECTED_2634,
  SV2V_UNCONNECTED_2635,SV2V_UNCONNECTED_2636,SV2V_UNCONNECTED_2637,
  SV2V_UNCONNECTED_2638,SV2V_UNCONNECTED_2639,SV2V_UNCONNECTED_2640,
  SV2V_UNCONNECTED_2641,SV2V_UNCONNECTED_2642,SV2V_UNCONNECTED_2643,
  SV2V_UNCONNECTED_2644,SV2V_UNCONNECTED_2645,SV2V_UNCONNECTED_2646,
  SV2V_UNCONNECTED_2647,SV2V_UNCONNECTED_2648,SV2V_UNCONNECTED_2649,
  SV2V_UNCONNECTED_2650,SV2V_UNCONNECTED_2651,SV2V_UNCONNECTED_2652,
  SV2V_UNCONNECTED_2653,SV2V_UNCONNECTED_2654,SV2V_UNCONNECTED_2655,
  SV2V_UNCONNECTED_2656,SV2V_UNCONNECTED_2657,SV2V_UNCONNECTED_2658,
  SV2V_UNCONNECTED_2659,SV2V_UNCONNECTED_2660,SV2V_UNCONNECTED_2661,
  SV2V_UNCONNECTED_2662,SV2V_UNCONNECTED_2663,SV2V_UNCONNECTED_2664,
  SV2V_UNCONNECTED_2665,SV2V_UNCONNECTED_2666,SV2V_UNCONNECTED_2667,SV2V_UNCONNECTED_2668,
  SV2V_UNCONNECTED_2669,SV2V_UNCONNECTED_2670,SV2V_UNCONNECTED_2671,
  SV2V_UNCONNECTED_2672,SV2V_UNCONNECTED_2673,SV2V_UNCONNECTED_2674,
  SV2V_UNCONNECTED_2675,SV2V_UNCONNECTED_2676,SV2V_UNCONNECTED_2677,
  SV2V_UNCONNECTED_2678,SV2V_UNCONNECTED_2679,SV2V_UNCONNECTED_2680,
  SV2V_UNCONNECTED_2681,SV2V_UNCONNECTED_2682,SV2V_UNCONNECTED_2683,
  SV2V_UNCONNECTED_2684,SV2V_UNCONNECTED_2685,SV2V_UNCONNECTED_2686,
  SV2V_UNCONNECTED_2687,SV2V_UNCONNECTED_2688,SV2V_UNCONNECTED_2689,
  SV2V_UNCONNECTED_2690,SV2V_UNCONNECTED_2691,SV2V_UNCONNECTED_2692,
  SV2V_UNCONNECTED_2693,SV2V_UNCONNECTED_2694,SV2V_UNCONNECTED_2695,
  SV2V_UNCONNECTED_2696,SV2V_UNCONNECTED_2697,SV2V_UNCONNECTED_2698,
  SV2V_UNCONNECTED_2699,SV2V_UNCONNECTED_2700,SV2V_UNCONNECTED_2701,
  SV2V_UNCONNECTED_2702,SV2V_UNCONNECTED_2703,SV2V_UNCONNECTED_2704,
  SV2V_UNCONNECTED_2705,SV2V_UNCONNECTED_2706,SV2V_UNCONNECTED_2707,SV2V_UNCONNECTED_2708,
  SV2V_UNCONNECTED_2709,SV2V_UNCONNECTED_2710,SV2V_UNCONNECTED_2711,
  SV2V_UNCONNECTED_2712,SV2V_UNCONNECTED_2713,SV2V_UNCONNECTED_2714,
  SV2V_UNCONNECTED_2715,SV2V_UNCONNECTED_2716,SV2V_UNCONNECTED_2717,
  SV2V_UNCONNECTED_2718,SV2V_UNCONNECTED_2719,SV2V_UNCONNECTED_2720,
  SV2V_UNCONNECTED_2721,SV2V_UNCONNECTED_2722,SV2V_UNCONNECTED_2723,
  SV2V_UNCONNECTED_2724,SV2V_UNCONNECTED_2725,SV2V_UNCONNECTED_2726,
  SV2V_UNCONNECTED_2727,SV2V_UNCONNECTED_2728,SV2V_UNCONNECTED_2729,
  SV2V_UNCONNECTED_2730,SV2V_UNCONNECTED_2731,SV2V_UNCONNECTED_2732,
  SV2V_UNCONNECTED_2733,SV2V_UNCONNECTED_2734,SV2V_UNCONNECTED_2735,
  SV2V_UNCONNECTED_2736,SV2V_UNCONNECTED_2737,SV2V_UNCONNECTED_2738,
  SV2V_UNCONNECTED_2739,SV2V_UNCONNECTED_2740,SV2V_UNCONNECTED_2741,
  SV2V_UNCONNECTED_2742,SV2V_UNCONNECTED_2743,SV2V_UNCONNECTED_2744,
  SV2V_UNCONNECTED_2745,SV2V_UNCONNECTED_2746,SV2V_UNCONNECTED_2747,SV2V_UNCONNECTED_2748,
  SV2V_UNCONNECTED_2749,SV2V_UNCONNECTED_2750,SV2V_UNCONNECTED_2751,
  SV2V_UNCONNECTED_2752,SV2V_UNCONNECTED_2753,SV2V_UNCONNECTED_2754,
  SV2V_UNCONNECTED_2755,SV2V_UNCONNECTED_2756,SV2V_UNCONNECTED_2757,
  SV2V_UNCONNECTED_2758,SV2V_UNCONNECTED_2759,SV2V_UNCONNECTED_2760,
  SV2V_UNCONNECTED_2761,SV2V_UNCONNECTED_2762,SV2V_UNCONNECTED_2763,
  SV2V_UNCONNECTED_2764,SV2V_UNCONNECTED_2765,SV2V_UNCONNECTED_2766,
  SV2V_UNCONNECTED_2767,SV2V_UNCONNECTED_2768,SV2V_UNCONNECTED_2769,
  SV2V_UNCONNECTED_2770,SV2V_UNCONNECTED_2771,SV2V_UNCONNECTED_2772,
  SV2V_UNCONNECTED_2773,SV2V_UNCONNECTED_2774,SV2V_UNCONNECTED_2775,
  SV2V_UNCONNECTED_2776,SV2V_UNCONNECTED_2777,SV2V_UNCONNECTED_2778,
  SV2V_UNCONNECTED_2779,SV2V_UNCONNECTED_2780,SV2V_UNCONNECTED_2781,
  SV2V_UNCONNECTED_2782,SV2V_UNCONNECTED_2783,SV2V_UNCONNECTED_2784,
  SV2V_UNCONNECTED_2785,SV2V_UNCONNECTED_2786,SV2V_UNCONNECTED_2787,SV2V_UNCONNECTED_2788,
  SV2V_UNCONNECTED_2789,SV2V_UNCONNECTED_2790,SV2V_UNCONNECTED_2791,
  SV2V_UNCONNECTED_2792,SV2V_UNCONNECTED_2793,SV2V_UNCONNECTED_2794,
  SV2V_UNCONNECTED_2795,SV2V_UNCONNECTED_2796,SV2V_UNCONNECTED_2797,
  SV2V_UNCONNECTED_2798,SV2V_UNCONNECTED_2799,SV2V_UNCONNECTED_2800,
  SV2V_UNCONNECTED_2801,SV2V_UNCONNECTED_2802,SV2V_UNCONNECTED_2803,
  SV2V_UNCONNECTED_2804,SV2V_UNCONNECTED_2805,SV2V_UNCONNECTED_2806,
  SV2V_UNCONNECTED_2807,SV2V_UNCONNECTED_2808,SV2V_UNCONNECTED_2809,
  SV2V_UNCONNECTED_2810,SV2V_UNCONNECTED_2811,SV2V_UNCONNECTED_2812,
  SV2V_UNCONNECTED_2813,SV2V_UNCONNECTED_2814,SV2V_UNCONNECTED_2815,
  SV2V_UNCONNECTED_2816,SV2V_UNCONNECTED_2817,SV2V_UNCONNECTED_2818,
  SV2V_UNCONNECTED_2819,SV2V_UNCONNECTED_2820,SV2V_UNCONNECTED_2821,
  SV2V_UNCONNECTED_2822,SV2V_UNCONNECTED_2823,SV2V_UNCONNECTED_2824,
  SV2V_UNCONNECTED_2825,SV2V_UNCONNECTED_2826,SV2V_UNCONNECTED_2827,SV2V_UNCONNECTED_2828,
  SV2V_UNCONNECTED_2829,SV2V_UNCONNECTED_2830,SV2V_UNCONNECTED_2831,
  SV2V_UNCONNECTED_2832,SV2V_UNCONNECTED_2833,SV2V_UNCONNECTED_2834,
  SV2V_UNCONNECTED_2835,SV2V_UNCONNECTED_2836,SV2V_UNCONNECTED_2837,
  SV2V_UNCONNECTED_2838,SV2V_UNCONNECTED_2839,SV2V_UNCONNECTED_2840,
  SV2V_UNCONNECTED_2841,SV2V_UNCONNECTED_2842,SV2V_UNCONNECTED_2843,
  SV2V_UNCONNECTED_2844,SV2V_UNCONNECTED_2845,SV2V_UNCONNECTED_2846,
  SV2V_UNCONNECTED_2847,SV2V_UNCONNECTED_2848,SV2V_UNCONNECTED_2849,
  SV2V_UNCONNECTED_2850,SV2V_UNCONNECTED_2851,SV2V_UNCONNECTED_2852,
  SV2V_UNCONNECTED_2853,SV2V_UNCONNECTED_2854,SV2V_UNCONNECTED_2855,
  SV2V_UNCONNECTED_2856,SV2V_UNCONNECTED_2857,SV2V_UNCONNECTED_2858,
  SV2V_UNCONNECTED_2859,SV2V_UNCONNECTED_2860,SV2V_UNCONNECTED_2861,
  SV2V_UNCONNECTED_2862,SV2V_UNCONNECTED_2863,SV2V_UNCONNECTED_2864,
  SV2V_UNCONNECTED_2865,SV2V_UNCONNECTED_2866,SV2V_UNCONNECTED_2867,SV2V_UNCONNECTED_2868,
  SV2V_UNCONNECTED_2869,SV2V_UNCONNECTED_2870,SV2V_UNCONNECTED_2871,
  SV2V_UNCONNECTED_2872,SV2V_UNCONNECTED_2873,SV2V_UNCONNECTED_2874,
  SV2V_UNCONNECTED_2875,SV2V_UNCONNECTED_2876,SV2V_UNCONNECTED_2877,
  SV2V_UNCONNECTED_2878,SV2V_UNCONNECTED_2879,SV2V_UNCONNECTED_2880,
  SV2V_UNCONNECTED_2881,SV2V_UNCONNECTED_2882,SV2V_UNCONNECTED_2883,
  SV2V_UNCONNECTED_2884,SV2V_UNCONNECTED_2885,SV2V_UNCONNECTED_2886,
  SV2V_UNCONNECTED_2887,SV2V_UNCONNECTED_2888,SV2V_UNCONNECTED_2889,
  SV2V_UNCONNECTED_2890,SV2V_UNCONNECTED_2891,SV2V_UNCONNECTED_2892,
  SV2V_UNCONNECTED_2893,SV2V_UNCONNECTED_2894,SV2V_UNCONNECTED_2895,
  SV2V_UNCONNECTED_2896,SV2V_UNCONNECTED_2897,SV2V_UNCONNECTED_2898,
  SV2V_UNCONNECTED_2899,SV2V_UNCONNECTED_2900,SV2V_UNCONNECTED_2901,
  SV2V_UNCONNECTED_2902,SV2V_UNCONNECTED_2903,SV2V_UNCONNECTED_2904,
  SV2V_UNCONNECTED_2905,SV2V_UNCONNECTED_2906,SV2V_UNCONNECTED_2907,SV2V_UNCONNECTED_2908,
  SV2V_UNCONNECTED_2909,SV2V_UNCONNECTED_2910,SV2V_UNCONNECTED_2911,
  SV2V_UNCONNECTED_2912,SV2V_UNCONNECTED_2913,SV2V_UNCONNECTED_2914,
  SV2V_UNCONNECTED_2915,SV2V_UNCONNECTED_2916,SV2V_UNCONNECTED_2917,
  SV2V_UNCONNECTED_2918,SV2V_UNCONNECTED_2919,SV2V_UNCONNECTED_2920,
  SV2V_UNCONNECTED_2921,SV2V_UNCONNECTED_2922,SV2V_UNCONNECTED_2923,
  SV2V_UNCONNECTED_2924,SV2V_UNCONNECTED_2925,SV2V_UNCONNECTED_2926,
  SV2V_UNCONNECTED_2927,SV2V_UNCONNECTED_2928,SV2V_UNCONNECTED_2929,
  SV2V_UNCONNECTED_2930,SV2V_UNCONNECTED_2931,SV2V_UNCONNECTED_2932,
  SV2V_UNCONNECTED_2933,SV2V_UNCONNECTED_2934,SV2V_UNCONNECTED_2935,
  SV2V_UNCONNECTED_2936,SV2V_UNCONNECTED_2937,SV2V_UNCONNECTED_2938,
  SV2V_UNCONNECTED_2939,SV2V_UNCONNECTED_2940,SV2V_UNCONNECTED_2941,
  SV2V_UNCONNECTED_2942,SV2V_UNCONNECTED_2943,SV2V_UNCONNECTED_2944,
  SV2V_UNCONNECTED_2945,SV2V_UNCONNECTED_2946,SV2V_UNCONNECTED_2947,SV2V_UNCONNECTED_2948,
  SV2V_UNCONNECTED_2949,SV2V_UNCONNECTED_2950,SV2V_UNCONNECTED_2951,
  SV2V_UNCONNECTED_2952,SV2V_UNCONNECTED_2953,SV2V_UNCONNECTED_2954,
  SV2V_UNCONNECTED_2955,SV2V_UNCONNECTED_2956,SV2V_UNCONNECTED_2957,
  SV2V_UNCONNECTED_2958,SV2V_UNCONNECTED_2959,SV2V_UNCONNECTED_2960,
  SV2V_UNCONNECTED_2961,SV2V_UNCONNECTED_2962,SV2V_UNCONNECTED_2963,
  SV2V_UNCONNECTED_2964,SV2V_UNCONNECTED_2965,SV2V_UNCONNECTED_2966,
  SV2V_UNCONNECTED_2967,SV2V_UNCONNECTED_2968,SV2V_UNCONNECTED_2969,
  SV2V_UNCONNECTED_2970,SV2V_UNCONNECTED_2971,SV2V_UNCONNECTED_2972,
  SV2V_UNCONNECTED_2973,SV2V_UNCONNECTED_2974,SV2V_UNCONNECTED_2975,
  SV2V_UNCONNECTED_2976,SV2V_UNCONNECTED_2977,SV2V_UNCONNECTED_2978,
  SV2V_UNCONNECTED_2979,SV2V_UNCONNECTED_2980,SV2V_UNCONNECTED_2981,
  SV2V_UNCONNECTED_2982,SV2V_UNCONNECTED_2983,SV2V_UNCONNECTED_2984,
  SV2V_UNCONNECTED_2985,SV2V_UNCONNECTED_2986,SV2V_UNCONNECTED_2987,SV2V_UNCONNECTED_2988,
  SV2V_UNCONNECTED_2989,SV2V_UNCONNECTED_2990,SV2V_UNCONNECTED_2991,
  SV2V_UNCONNECTED_2992,SV2V_UNCONNECTED_2993,SV2V_UNCONNECTED_2994,
  SV2V_UNCONNECTED_2995,SV2V_UNCONNECTED_2996,SV2V_UNCONNECTED_2997,
  SV2V_UNCONNECTED_2998,SV2V_UNCONNECTED_2999,SV2V_UNCONNECTED_3000,
  SV2V_UNCONNECTED_3001,SV2V_UNCONNECTED_3002,SV2V_UNCONNECTED_3003,
  SV2V_UNCONNECTED_3004,SV2V_UNCONNECTED_3005,SV2V_UNCONNECTED_3006,
  SV2V_UNCONNECTED_3007,SV2V_UNCONNECTED_3008,SV2V_UNCONNECTED_3009,
  SV2V_UNCONNECTED_3010,SV2V_UNCONNECTED_3011,SV2V_UNCONNECTED_3012,
  SV2V_UNCONNECTED_3013,SV2V_UNCONNECTED_3014,SV2V_UNCONNECTED_3015,
  SV2V_UNCONNECTED_3016,SV2V_UNCONNECTED_3017,SV2V_UNCONNECTED_3018,
  SV2V_UNCONNECTED_3019,SV2V_UNCONNECTED_3020,SV2V_UNCONNECTED_3021,
  SV2V_UNCONNECTED_3022,SV2V_UNCONNECTED_3023,SV2V_UNCONNECTED_3024,
  SV2V_UNCONNECTED_3025,SV2V_UNCONNECTED_3026,SV2V_UNCONNECTED_3027,SV2V_UNCONNECTED_3028,
  SV2V_UNCONNECTED_3029,SV2V_UNCONNECTED_3030,SV2V_UNCONNECTED_3031,
  SV2V_UNCONNECTED_3032,SV2V_UNCONNECTED_3033,SV2V_UNCONNECTED_3034,
  SV2V_UNCONNECTED_3035,SV2V_UNCONNECTED_3036,SV2V_UNCONNECTED_3037,
  SV2V_UNCONNECTED_3038,SV2V_UNCONNECTED_3039,SV2V_UNCONNECTED_3040,
  SV2V_UNCONNECTED_3041,SV2V_UNCONNECTED_3042,SV2V_UNCONNECTED_3043,
  SV2V_UNCONNECTED_3044,SV2V_UNCONNECTED_3045,SV2V_UNCONNECTED_3046,
  SV2V_UNCONNECTED_3047,SV2V_UNCONNECTED_3048,SV2V_UNCONNECTED_3049,
  SV2V_UNCONNECTED_3050,SV2V_UNCONNECTED_3051,SV2V_UNCONNECTED_3052,
  SV2V_UNCONNECTED_3053,SV2V_UNCONNECTED_3054,SV2V_UNCONNECTED_3055,
  SV2V_UNCONNECTED_3056,SV2V_UNCONNECTED_3057,SV2V_UNCONNECTED_3058,
  SV2V_UNCONNECTED_3059,SV2V_UNCONNECTED_3060,SV2V_UNCONNECTED_3061,
  SV2V_UNCONNECTED_3062,SV2V_UNCONNECTED_3063,SV2V_UNCONNECTED_3064,
  SV2V_UNCONNECTED_3065,SV2V_UNCONNECTED_3066,SV2V_UNCONNECTED_3067,SV2V_UNCONNECTED_3068,
  SV2V_UNCONNECTED_3069,SV2V_UNCONNECTED_3070,SV2V_UNCONNECTED_3071,
  SV2V_UNCONNECTED_3072,SV2V_UNCONNECTED_3073,SV2V_UNCONNECTED_3074,
  SV2V_UNCONNECTED_3075,SV2V_UNCONNECTED_3076,SV2V_UNCONNECTED_3077,
  SV2V_UNCONNECTED_3078,SV2V_UNCONNECTED_3079,SV2V_UNCONNECTED_3080,
  SV2V_UNCONNECTED_3081,SV2V_UNCONNECTED_3082,SV2V_UNCONNECTED_3083,
  SV2V_UNCONNECTED_3084,SV2V_UNCONNECTED_3085,SV2V_UNCONNECTED_3086,
  SV2V_UNCONNECTED_3087,SV2V_UNCONNECTED_3088,SV2V_UNCONNECTED_3089,
  SV2V_UNCONNECTED_3090,SV2V_UNCONNECTED_3091,SV2V_UNCONNECTED_3092,
  SV2V_UNCONNECTED_3093,SV2V_UNCONNECTED_3094,SV2V_UNCONNECTED_3095,
  SV2V_UNCONNECTED_3096,SV2V_UNCONNECTED_3097,SV2V_UNCONNECTED_3098,
  SV2V_UNCONNECTED_3099,SV2V_UNCONNECTED_3100,SV2V_UNCONNECTED_3101,
  SV2V_UNCONNECTED_3102,SV2V_UNCONNECTED_3103,SV2V_UNCONNECTED_3104,
  SV2V_UNCONNECTED_3105,SV2V_UNCONNECTED_3106,SV2V_UNCONNECTED_3107,SV2V_UNCONNECTED_3108,
  SV2V_UNCONNECTED_3109,SV2V_UNCONNECTED_3110,SV2V_UNCONNECTED_3111,
  SV2V_UNCONNECTED_3112,SV2V_UNCONNECTED_3113,SV2V_UNCONNECTED_3114,
  SV2V_UNCONNECTED_3115,SV2V_UNCONNECTED_3116,SV2V_UNCONNECTED_3117,
  SV2V_UNCONNECTED_3118,SV2V_UNCONNECTED_3119,SV2V_UNCONNECTED_3120,
  SV2V_UNCONNECTED_3121,SV2V_UNCONNECTED_3122,SV2V_UNCONNECTED_3123,
  SV2V_UNCONNECTED_3124,SV2V_UNCONNECTED_3125,SV2V_UNCONNECTED_3126,
  SV2V_UNCONNECTED_3127,SV2V_UNCONNECTED_3128,SV2V_UNCONNECTED_3129,
  SV2V_UNCONNECTED_3130,SV2V_UNCONNECTED_3131,SV2V_UNCONNECTED_3132,
  SV2V_UNCONNECTED_3133,SV2V_UNCONNECTED_3134,SV2V_UNCONNECTED_3135,
  SV2V_UNCONNECTED_3136,SV2V_UNCONNECTED_3137,SV2V_UNCONNECTED_3138,
  SV2V_UNCONNECTED_3139,SV2V_UNCONNECTED_3140,SV2V_UNCONNECTED_3141,
  SV2V_UNCONNECTED_3142,SV2V_UNCONNECTED_3143,SV2V_UNCONNECTED_3144,
  SV2V_UNCONNECTED_3145,SV2V_UNCONNECTED_3146,SV2V_UNCONNECTED_3147,SV2V_UNCONNECTED_3148,
  SV2V_UNCONNECTED_3149,SV2V_UNCONNECTED_3150,SV2V_UNCONNECTED_3151,
  SV2V_UNCONNECTED_3152,SV2V_UNCONNECTED_3153,SV2V_UNCONNECTED_3154,
  SV2V_UNCONNECTED_3155,SV2V_UNCONNECTED_3156,SV2V_UNCONNECTED_3157,
  SV2V_UNCONNECTED_3158,SV2V_UNCONNECTED_3159,SV2V_UNCONNECTED_3160,
  SV2V_UNCONNECTED_3161,SV2V_UNCONNECTED_3162,SV2V_UNCONNECTED_3163,
  SV2V_UNCONNECTED_3164,SV2V_UNCONNECTED_3165,SV2V_UNCONNECTED_3166,
  SV2V_UNCONNECTED_3167,SV2V_UNCONNECTED_3168,SV2V_UNCONNECTED_3169,
  SV2V_UNCONNECTED_3170,SV2V_UNCONNECTED_3171,SV2V_UNCONNECTED_3172,
  SV2V_UNCONNECTED_3173,SV2V_UNCONNECTED_3174,SV2V_UNCONNECTED_3175,
  SV2V_UNCONNECTED_3176,SV2V_UNCONNECTED_3177,SV2V_UNCONNECTED_3178,
  SV2V_UNCONNECTED_3179,SV2V_UNCONNECTED_3180,SV2V_UNCONNECTED_3181,
  SV2V_UNCONNECTED_3182,SV2V_UNCONNECTED_3183,SV2V_UNCONNECTED_3184,
  SV2V_UNCONNECTED_3185,SV2V_UNCONNECTED_3186,SV2V_UNCONNECTED_3187,SV2V_UNCONNECTED_3188,
  SV2V_UNCONNECTED_3189,SV2V_UNCONNECTED_3190,SV2V_UNCONNECTED_3191,
  SV2V_UNCONNECTED_3192,SV2V_UNCONNECTED_3193,SV2V_UNCONNECTED_3194,
  SV2V_UNCONNECTED_3195,SV2V_UNCONNECTED_3196,SV2V_UNCONNECTED_3197,
  SV2V_UNCONNECTED_3198,SV2V_UNCONNECTED_3199,SV2V_UNCONNECTED_3200,
  SV2V_UNCONNECTED_3201,SV2V_UNCONNECTED_3202,SV2V_UNCONNECTED_3203,
  SV2V_UNCONNECTED_3204,SV2V_UNCONNECTED_3205,SV2V_UNCONNECTED_3206,
  SV2V_UNCONNECTED_3207,SV2V_UNCONNECTED_3208,SV2V_UNCONNECTED_3209,
  SV2V_UNCONNECTED_3210,SV2V_UNCONNECTED_3211,SV2V_UNCONNECTED_3212,
  SV2V_UNCONNECTED_3213,SV2V_UNCONNECTED_3214,SV2V_UNCONNECTED_3215,
  SV2V_UNCONNECTED_3216,SV2V_UNCONNECTED_3217,SV2V_UNCONNECTED_3218,
  SV2V_UNCONNECTED_3219,SV2V_UNCONNECTED_3220,SV2V_UNCONNECTED_3221,
  SV2V_UNCONNECTED_3222,SV2V_UNCONNECTED_3223,SV2V_UNCONNECTED_3224,
  SV2V_UNCONNECTED_3225,SV2V_UNCONNECTED_3226,SV2V_UNCONNECTED_3227,SV2V_UNCONNECTED_3228,
  SV2V_UNCONNECTED_3229,SV2V_UNCONNECTED_3230,SV2V_UNCONNECTED_3231,
  SV2V_UNCONNECTED_3232,SV2V_UNCONNECTED_3233,SV2V_UNCONNECTED_3234,
  SV2V_UNCONNECTED_3235,SV2V_UNCONNECTED_3236,SV2V_UNCONNECTED_3237,
  SV2V_UNCONNECTED_3238,SV2V_UNCONNECTED_3239,SV2V_UNCONNECTED_3240,
  SV2V_UNCONNECTED_3241,SV2V_UNCONNECTED_3242,SV2V_UNCONNECTED_3243,
  SV2V_UNCONNECTED_3244,SV2V_UNCONNECTED_3245,SV2V_UNCONNECTED_3246,
  SV2V_UNCONNECTED_3247,SV2V_UNCONNECTED_3248,SV2V_UNCONNECTED_3249,
  SV2V_UNCONNECTED_3250,SV2V_UNCONNECTED_3251,SV2V_UNCONNECTED_3252,
  SV2V_UNCONNECTED_3253,SV2V_UNCONNECTED_3254,SV2V_UNCONNECTED_3255,
  SV2V_UNCONNECTED_3256,SV2V_UNCONNECTED_3257,SV2V_UNCONNECTED_3258,
  SV2V_UNCONNECTED_3259,SV2V_UNCONNECTED_3260,SV2V_UNCONNECTED_3261,
  SV2V_UNCONNECTED_3262,SV2V_UNCONNECTED_3263,SV2V_UNCONNECTED_3264,
  SV2V_UNCONNECTED_3265,SV2V_UNCONNECTED_3266,SV2V_UNCONNECTED_3267,SV2V_UNCONNECTED_3268,
  SV2V_UNCONNECTED_3269,SV2V_UNCONNECTED_3270,SV2V_UNCONNECTED_3271,
  SV2V_UNCONNECTED_3272,SV2V_UNCONNECTED_3273,SV2V_UNCONNECTED_3274,
  SV2V_UNCONNECTED_3275,SV2V_UNCONNECTED_3276,SV2V_UNCONNECTED_3277,
  SV2V_UNCONNECTED_3278,SV2V_UNCONNECTED_3279,SV2V_UNCONNECTED_3280,
  SV2V_UNCONNECTED_3281,SV2V_UNCONNECTED_3282,SV2V_UNCONNECTED_3283,
  SV2V_UNCONNECTED_3284,SV2V_UNCONNECTED_3285,SV2V_UNCONNECTED_3286,
  SV2V_UNCONNECTED_3287,SV2V_UNCONNECTED_3288,SV2V_UNCONNECTED_3289,
  SV2V_UNCONNECTED_3290,SV2V_UNCONNECTED_3291,SV2V_UNCONNECTED_3292,
  SV2V_UNCONNECTED_3293,SV2V_UNCONNECTED_3294,SV2V_UNCONNECTED_3295,
  SV2V_UNCONNECTED_3296,SV2V_UNCONNECTED_3297,SV2V_UNCONNECTED_3298,
  SV2V_UNCONNECTED_3299,SV2V_UNCONNECTED_3300,SV2V_UNCONNECTED_3301,
  SV2V_UNCONNECTED_3302,SV2V_UNCONNECTED_3303,SV2V_UNCONNECTED_3304,
  SV2V_UNCONNECTED_3305,SV2V_UNCONNECTED_3306,SV2V_UNCONNECTED_3307,SV2V_UNCONNECTED_3308,
  SV2V_UNCONNECTED_3309,SV2V_UNCONNECTED_3310,SV2V_UNCONNECTED_3311,
  SV2V_UNCONNECTED_3312,SV2V_UNCONNECTED_3313,SV2V_UNCONNECTED_3314,
  SV2V_UNCONNECTED_3315,SV2V_UNCONNECTED_3316,SV2V_UNCONNECTED_3317,
  SV2V_UNCONNECTED_3318,SV2V_UNCONNECTED_3319,SV2V_UNCONNECTED_3320,
  SV2V_UNCONNECTED_3321,SV2V_UNCONNECTED_3322,SV2V_UNCONNECTED_3323,
  SV2V_UNCONNECTED_3324,SV2V_UNCONNECTED_3325,SV2V_UNCONNECTED_3326,
  SV2V_UNCONNECTED_3327,SV2V_UNCONNECTED_3328,SV2V_UNCONNECTED_3329,
  SV2V_UNCONNECTED_3330,SV2V_UNCONNECTED_3331,SV2V_UNCONNECTED_3332,
  SV2V_UNCONNECTED_3333,SV2V_UNCONNECTED_3334,SV2V_UNCONNECTED_3335,
  SV2V_UNCONNECTED_3336,SV2V_UNCONNECTED_3337,SV2V_UNCONNECTED_3338,
  SV2V_UNCONNECTED_3339,SV2V_UNCONNECTED_3340,SV2V_UNCONNECTED_3341,
  SV2V_UNCONNECTED_3342,SV2V_UNCONNECTED_3343,SV2V_UNCONNECTED_3344,
  SV2V_UNCONNECTED_3345,SV2V_UNCONNECTED_3346,SV2V_UNCONNECTED_3347,SV2V_UNCONNECTED_3348,
  SV2V_UNCONNECTED_3349,SV2V_UNCONNECTED_3350,SV2V_UNCONNECTED_3351,
  SV2V_UNCONNECTED_3352,SV2V_UNCONNECTED_3353,SV2V_UNCONNECTED_3354,
  SV2V_UNCONNECTED_3355,SV2V_UNCONNECTED_3356,SV2V_UNCONNECTED_3357,
  SV2V_UNCONNECTED_3358,SV2V_UNCONNECTED_3359,SV2V_UNCONNECTED_3360,
  SV2V_UNCONNECTED_3361,SV2V_UNCONNECTED_3362,SV2V_UNCONNECTED_3363,
  SV2V_UNCONNECTED_3364,SV2V_UNCONNECTED_3365,SV2V_UNCONNECTED_3366,
  SV2V_UNCONNECTED_3367,SV2V_UNCONNECTED_3368,SV2V_UNCONNECTED_3369,
  SV2V_UNCONNECTED_3370,SV2V_UNCONNECTED_3371,SV2V_UNCONNECTED_3372,
  SV2V_UNCONNECTED_3373,SV2V_UNCONNECTED_3374,SV2V_UNCONNECTED_3375,
  SV2V_UNCONNECTED_3376,SV2V_UNCONNECTED_3377,SV2V_UNCONNECTED_3378,
  SV2V_UNCONNECTED_3379,SV2V_UNCONNECTED_3380,SV2V_UNCONNECTED_3381,
  SV2V_UNCONNECTED_3382,SV2V_UNCONNECTED_3383,SV2V_UNCONNECTED_3384,
  SV2V_UNCONNECTED_3385,SV2V_UNCONNECTED_3386,SV2V_UNCONNECTED_3387,SV2V_UNCONNECTED_3388,
  SV2V_UNCONNECTED_3389,SV2V_UNCONNECTED_3390,SV2V_UNCONNECTED_3391,
  SV2V_UNCONNECTED_3392,SV2V_UNCONNECTED_3393,SV2V_UNCONNECTED_3394,
  SV2V_UNCONNECTED_3395,SV2V_UNCONNECTED_3396,SV2V_UNCONNECTED_3397,
  SV2V_UNCONNECTED_3398,SV2V_UNCONNECTED_3399,SV2V_UNCONNECTED_3400,
  SV2V_UNCONNECTED_3401,SV2V_UNCONNECTED_3402,SV2V_UNCONNECTED_3403,
  SV2V_UNCONNECTED_3404,SV2V_UNCONNECTED_3405,SV2V_UNCONNECTED_3406,
  SV2V_UNCONNECTED_3407,SV2V_UNCONNECTED_3408,SV2V_UNCONNECTED_3409,
  SV2V_UNCONNECTED_3410,SV2V_UNCONNECTED_3411,SV2V_UNCONNECTED_3412,
  SV2V_UNCONNECTED_3413,SV2V_UNCONNECTED_3414,SV2V_UNCONNECTED_3415,
  SV2V_UNCONNECTED_3416,SV2V_UNCONNECTED_3417,SV2V_UNCONNECTED_3418,
  SV2V_UNCONNECTED_3419,SV2V_UNCONNECTED_3420,SV2V_UNCONNECTED_3421,
  SV2V_UNCONNECTED_3422,SV2V_UNCONNECTED_3423,SV2V_UNCONNECTED_3424,
  SV2V_UNCONNECTED_3425,SV2V_UNCONNECTED_3426,SV2V_UNCONNECTED_3427,SV2V_UNCONNECTED_3428,
  SV2V_UNCONNECTED_3429,SV2V_UNCONNECTED_3430,SV2V_UNCONNECTED_3431,
  SV2V_UNCONNECTED_3432,SV2V_UNCONNECTED_3433,SV2V_UNCONNECTED_3434,
  SV2V_UNCONNECTED_3435,SV2V_UNCONNECTED_3436,SV2V_UNCONNECTED_3437,
  SV2V_UNCONNECTED_3438,SV2V_UNCONNECTED_3439,SV2V_UNCONNECTED_3440,
  SV2V_UNCONNECTED_3441,SV2V_UNCONNECTED_3442,SV2V_UNCONNECTED_3443,
  SV2V_UNCONNECTED_3444,SV2V_UNCONNECTED_3445,SV2V_UNCONNECTED_3446,
  SV2V_UNCONNECTED_3447,SV2V_UNCONNECTED_3448,SV2V_UNCONNECTED_3449,
  SV2V_UNCONNECTED_3450,SV2V_UNCONNECTED_3451,SV2V_UNCONNECTED_3452,
  SV2V_UNCONNECTED_3453,SV2V_UNCONNECTED_3454,SV2V_UNCONNECTED_3455,
  SV2V_UNCONNECTED_3456,SV2V_UNCONNECTED_3457,SV2V_UNCONNECTED_3458,
  SV2V_UNCONNECTED_3459,SV2V_UNCONNECTED_3460,SV2V_UNCONNECTED_3461,
  SV2V_UNCONNECTED_3462,SV2V_UNCONNECTED_3463,SV2V_UNCONNECTED_3464,
  SV2V_UNCONNECTED_3465,SV2V_UNCONNECTED_3466,SV2V_UNCONNECTED_3467,SV2V_UNCONNECTED_3468,
  SV2V_UNCONNECTED_3469,SV2V_UNCONNECTED_3470,SV2V_UNCONNECTED_3471,
  SV2V_UNCONNECTED_3472,SV2V_UNCONNECTED_3473,SV2V_UNCONNECTED_3474,
  SV2V_UNCONNECTED_3475,SV2V_UNCONNECTED_3476,SV2V_UNCONNECTED_3477,
  SV2V_UNCONNECTED_3478,SV2V_UNCONNECTED_3479,SV2V_UNCONNECTED_3480,
  SV2V_UNCONNECTED_3481,SV2V_UNCONNECTED_3482,SV2V_UNCONNECTED_3483,
  SV2V_UNCONNECTED_3484,SV2V_UNCONNECTED_3485,SV2V_UNCONNECTED_3486,
  SV2V_UNCONNECTED_3487,SV2V_UNCONNECTED_3488,SV2V_UNCONNECTED_3489,
  SV2V_UNCONNECTED_3490,SV2V_UNCONNECTED_3491,SV2V_UNCONNECTED_3492,
  SV2V_UNCONNECTED_3493,SV2V_UNCONNECTED_3494,SV2V_UNCONNECTED_3495,
  SV2V_UNCONNECTED_3496,SV2V_UNCONNECTED_3497,SV2V_UNCONNECTED_3498,
  SV2V_UNCONNECTED_3499,SV2V_UNCONNECTED_3500,SV2V_UNCONNECTED_3501,
  SV2V_UNCONNECTED_3502,SV2V_UNCONNECTED_3503,SV2V_UNCONNECTED_3504,
  SV2V_UNCONNECTED_3505,SV2V_UNCONNECTED_3506,SV2V_UNCONNECTED_3507,SV2V_UNCONNECTED_3508,
  SV2V_UNCONNECTED_3509,SV2V_UNCONNECTED_3510,SV2V_UNCONNECTED_3511,
  SV2V_UNCONNECTED_3512,SV2V_UNCONNECTED_3513,SV2V_UNCONNECTED_3514,
  SV2V_UNCONNECTED_3515,SV2V_UNCONNECTED_3516,SV2V_UNCONNECTED_3517,
  SV2V_UNCONNECTED_3518,SV2V_UNCONNECTED_3519,SV2V_UNCONNECTED_3520,
  SV2V_UNCONNECTED_3521,SV2V_UNCONNECTED_3522,SV2V_UNCONNECTED_3523,
  SV2V_UNCONNECTED_3524,SV2V_UNCONNECTED_3525,SV2V_UNCONNECTED_3526,
  SV2V_UNCONNECTED_3527,SV2V_UNCONNECTED_3528,SV2V_UNCONNECTED_3529,
  SV2V_UNCONNECTED_3530,SV2V_UNCONNECTED_3531,SV2V_UNCONNECTED_3532,
  SV2V_UNCONNECTED_3533,SV2V_UNCONNECTED_3534,SV2V_UNCONNECTED_3535,
  SV2V_UNCONNECTED_3536,SV2V_UNCONNECTED_3537,SV2V_UNCONNECTED_3538,
  SV2V_UNCONNECTED_3539,SV2V_UNCONNECTED_3540,SV2V_UNCONNECTED_3541,
  SV2V_UNCONNECTED_3542,SV2V_UNCONNECTED_3543,SV2V_UNCONNECTED_3544,
  SV2V_UNCONNECTED_3545,SV2V_UNCONNECTED_3546,SV2V_UNCONNECTED_3547,SV2V_UNCONNECTED_3548,
  SV2V_UNCONNECTED_3549,SV2V_UNCONNECTED_3550,SV2V_UNCONNECTED_3551,
  SV2V_UNCONNECTED_3552,SV2V_UNCONNECTED_3553,SV2V_UNCONNECTED_3554,
  SV2V_UNCONNECTED_3555,SV2V_UNCONNECTED_3556,SV2V_UNCONNECTED_3557,
  SV2V_UNCONNECTED_3558,SV2V_UNCONNECTED_3559,SV2V_UNCONNECTED_3560,
  SV2V_UNCONNECTED_3561,SV2V_UNCONNECTED_3562,SV2V_UNCONNECTED_3563,
  SV2V_UNCONNECTED_3564,SV2V_UNCONNECTED_3565,SV2V_UNCONNECTED_3566,
  SV2V_UNCONNECTED_3567,SV2V_UNCONNECTED_3568,SV2V_UNCONNECTED_3569,
  SV2V_UNCONNECTED_3570,SV2V_UNCONNECTED_3571,SV2V_UNCONNECTED_3572,
  SV2V_UNCONNECTED_3573,SV2V_UNCONNECTED_3574,SV2V_UNCONNECTED_3575,
  SV2V_UNCONNECTED_3576,SV2V_UNCONNECTED_3577,SV2V_UNCONNECTED_3578,
  SV2V_UNCONNECTED_3579,SV2V_UNCONNECTED_3580,SV2V_UNCONNECTED_3581,
  SV2V_UNCONNECTED_3582,SV2V_UNCONNECTED_3583,SV2V_UNCONNECTED_3584,
  SV2V_UNCONNECTED_3585,SV2V_UNCONNECTED_3586,SV2V_UNCONNECTED_3587,SV2V_UNCONNECTED_3588,
  SV2V_UNCONNECTED_3589,SV2V_UNCONNECTED_3590,SV2V_UNCONNECTED_3591,
  SV2V_UNCONNECTED_3592,SV2V_UNCONNECTED_3593,SV2V_UNCONNECTED_3594,
  SV2V_UNCONNECTED_3595,SV2V_UNCONNECTED_3596,SV2V_UNCONNECTED_3597,
  SV2V_UNCONNECTED_3598,SV2V_UNCONNECTED_3599,SV2V_UNCONNECTED_3600,
  SV2V_UNCONNECTED_3601,SV2V_UNCONNECTED_3602,SV2V_UNCONNECTED_3603,
  SV2V_UNCONNECTED_3604,SV2V_UNCONNECTED_3605,SV2V_UNCONNECTED_3606,
  SV2V_UNCONNECTED_3607,SV2V_UNCONNECTED_3608,SV2V_UNCONNECTED_3609,
  SV2V_UNCONNECTED_3610,SV2V_UNCONNECTED_3611,SV2V_UNCONNECTED_3612,
  SV2V_UNCONNECTED_3613,SV2V_UNCONNECTED_3614,SV2V_UNCONNECTED_3615,
  SV2V_UNCONNECTED_3616,SV2V_UNCONNECTED_3617,SV2V_UNCONNECTED_3618,
  SV2V_UNCONNECTED_3619,SV2V_UNCONNECTED_3620,SV2V_UNCONNECTED_3621,
  SV2V_UNCONNECTED_3622,SV2V_UNCONNECTED_3623,SV2V_UNCONNECTED_3624,
  SV2V_UNCONNECTED_3625,SV2V_UNCONNECTED_3626,SV2V_UNCONNECTED_3627,SV2V_UNCONNECTED_3628,
  SV2V_UNCONNECTED_3629,SV2V_UNCONNECTED_3630,SV2V_UNCONNECTED_3631,
  SV2V_UNCONNECTED_3632,SV2V_UNCONNECTED_3633,SV2V_UNCONNECTED_3634,
  SV2V_UNCONNECTED_3635,SV2V_UNCONNECTED_3636,SV2V_UNCONNECTED_3637,
  SV2V_UNCONNECTED_3638,SV2V_UNCONNECTED_3639,SV2V_UNCONNECTED_3640,
  SV2V_UNCONNECTED_3641,SV2V_UNCONNECTED_3642,SV2V_UNCONNECTED_3643,
  SV2V_UNCONNECTED_3644,SV2V_UNCONNECTED_3645,SV2V_UNCONNECTED_3646,
  SV2V_UNCONNECTED_3647,SV2V_UNCONNECTED_3648,SV2V_UNCONNECTED_3649,
  SV2V_UNCONNECTED_3650,SV2V_UNCONNECTED_3651,SV2V_UNCONNECTED_3652,
  SV2V_UNCONNECTED_3653,SV2V_UNCONNECTED_3654,SV2V_UNCONNECTED_3655,
  SV2V_UNCONNECTED_3656,SV2V_UNCONNECTED_3657,SV2V_UNCONNECTED_3658,
  SV2V_UNCONNECTED_3659,SV2V_UNCONNECTED_3660,SV2V_UNCONNECTED_3661,
  SV2V_UNCONNECTED_3662,SV2V_UNCONNECTED_3663,SV2V_UNCONNECTED_3664,
  SV2V_UNCONNECTED_3665,SV2V_UNCONNECTED_3666,SV2V_UNCONNECTED_3667,SV2V_UNCONNECTED_3668,
  SV2V_UNCONNECTED_3669,SV2V_UNCONNECTED_3670,SV2V_UNCONNECTED_3671,
  SV2V_UNCONNECTED_3672,SV2V_UNCONNECTED_3673,SV2V_UNCONNECTED_3674,
  SV2V_UNCONNECTED_3675,SV2V_UNCONNECTED_3676,SV2V_UNCONNECTED_3677,
  SV2V_UNCONNECTED_3678,SV2V_UNCONNECTED_3679,SV2V_UNCONNECTED_3680,
  SV2V_UNCONNECTED_3681,SV2V_UNCONNECTED_3682,SV2V_UNCONNECTED_3683,
  SV2V_UNCONNECTED_3684,SV2V_UNCONNECTED_3685,SV2V_UNCONNECTED_3686,
  SV2V_UNCONNECTED_3687,SV2V_UNCONNECTED_3688,SV2V_UNCONNECTED_3689,
  SV2V_UNCONNECTED_3690,SV2V_UNCONNECTED_3691,SV2V_UNCONNECTED_3692,
  SV2V_UNCONNECTED_3693,SV2V_UNCONNECTED_3694,SV2V_UNCONNECTED_3695,
  SV2V_UNCONNECTED_3696,SV2V_UNCONNECTED_3697,SV2V_UNCONNECTED_3698,
  SV2V_UNCONNECTED_3699,SV2V_UNCONNECTED_3700,SV2V_UNCONNECTED_3701,
  SV2V_UNCONNECTED_3702,SV2V_UNCONNECTED_3703,SV2V_UNCONNECTED_3704,
  SV2V_UNCONNECTED_3705,SV2V_UNCONNECTED_3706,SV2V_UNCONNECTED_3707,SV2V_UNCONNECTED_3708,
  SV2V_UNCONNECTED_3709,SV2V_UNCONNECTED_3710,SV2V_UNCONNECTED_3711,
  SV2V_UNCONNECTED_3712,SV2V_UNCONNECTED_3713,SV2V_UNCONNECTED_3714,
  SV2V_UNCONNECTED_3715,SV2V_UNCONNECTED_3716,SV2V_UNCONNECTED_3717,
  SV2V_UNCONNECTED_3718,SV2V_UNCONNECTED_3719,SV2V_UNCONNECTED_3720,
  SV2V_UNCONNECTED_3721,SV2V_UNCONNECTED_3722,SV2V_UNCONNECTED_3723,
  SV2V_UNCONNECTED_3724,SV2V_UNCONNECTED_3725,SV2V_UNCONNECTED_3726,
  SV2V_UNCONNECTED_3727,SV2V_UNCONNECTED_3728,SV2V_UNCONNECTED_3729,
  SV2V_UNCONNECTED_3730,SV2V_UNCONNECTED_3731,SV2V_UNCONNECTED_3732,
  SV2V_UNCONNECTED_3733,SV2V_UNCONNECTED_3734,SV2V_UNCONNECTED_3735,
  SV2V_UNCONNECTED_3736,SV2V_UNCONNECTED_3737,SV2V_UNCONNECTED_3738,
  SV2V_UNCONNECTED_3739,SV2V_UNCONNECTED_3740,SV2V_UNCONNECTED_3741,
  SV2V_UNCONNECTED_3742,SV2V_UNCONNECTED_3743,SV2V_UNCONNECTED_3744,
  SV2V_UNCONNECTED_3745,SV2V_UNCONNECTED_3746,SV2V_UNCONNECTED_3747,SV2V_UNCONNECTED_3748,
  SV2V_UNCONNECTED_3749,SV2V_UNCONNECTED_3750,SV2V_UNCONNECTED_3751,
  SV2V_UNCONNECTED_3752,SV2V_UNCONNECTED_3753,SV2V_UNCONNECTED_3754,
  SV2V_UNCONNECTED_3755,SV2V_UNCONNECTED_3756,SV2V_UNCONNECTED_3757,
  SV2V_UNCONNECTED_3758,SV2V_UNCONNECTED_3759,SV2V_UNCONNECTED_3760,
  SV2V_UNCONNECTED_3761,SV2V_UNCONNECTED_3762,SV2V_UNCONNECTED_3763,
  SV2V_UNCONNECTED_3764,SV2V_UNCONNECTED_3765,SV2V_UNCONNECTED_3766,
  SV2V_UNCONNECTED_3767,SV2V_UNCONNECTED_3768,SV2V_UNCONNECTED_3769,
  SV2V_UNCONNECTED_3770,SV2V_UNCONNECTED_3771,SV2V_UNCONNECTED_3772,
  SV2V_UNCONNECTED_3773,SV2V_UNCONNECTED_3774,SV2V_UNCONNECTED_3775,
  SV2V_UNCONNECTED_3776,SV2V_UNCONNECTED_3777,SV2V_UNCONNECTED_3778,
  SV2V_UNCONNECTED_3779,SV2V_UNCONNECTED_3780,SV2V_UNCONNECTED_3781,
  SV2V_UNCONNECTED_3782,SV2V_UNCONNECTED_3783,SV2V_UNCONNECTED_3784,
  SV2V_UNCONNECTED_3785,SV2V_UNCONNECTED_3786,SV2V_UNCONNECTED_3787,SV2V_UNCONNECTED_3788,
  SV2V_UNCONNECTED_3789,SV2V_UNCONNECTED_3790,SV2V_UNCONNECTED_3791,
  SV2V_UNCONNECTED_3792,SV2V_UNCONNECTED_3793,SV2V_UNCONNECTED_3794,
  SV2V_UNCONNECTED_3795,SV2V_UNCONNECTED_3796,SV2V_UNCONNECTED_3797,
  SV2V_UNCONNECTED_3798,SV2V_UNCONNECTED_3799,SV2V_UNCONNECTED_3800,
  SV2V_UNCONNECTED_3801,SV2V_UNCONNECTED_3802,SV2V_UNCONNECTED_3803,
  SV2V_UNCONNECTED_3804,SV2V_UNCONNECTED_3805,SV2V_UNCONNECTED_3806,
  SV2V_UNCONNECTED_3807,SV2V_UNCONNECTED_3808,SV2V_UNCONNECTED_3809,
  SV2V_UNCONNECTED_3810,SV2V_UNCONNECTED_3811,SV2V_UNCONNECTED_3812,
  SV2V_UNCONNECTED_3813,SV2V_UNCONNECTED_3814,SV2V_UNCONNECTED_3815,
  SV2V_UNCONNECTED_3816,SV2V_UNCONNECTED_3817,SV2V_UNCONNECTED_3818,
  SV2V_UNCONNECTED_3819,SV2V_UNCONNECTED_3820,SV2V_UNCONNECTED_3821,
  SV2V_UNCONNECTED_3822,SV2V_UNCONNECTED_3823,SV2V_UNCONNECTED_3824,
  SV2V_UNCONNECTED_3825,SV2V_UNCONNECTED_3826,SV2V_UNCONNECTED_3827,SV2V_UNCONNECTED_3828,
  SV2V_UNCONNECTED_3829,SV2V_UNCONNECTED_3830,SV2V_UNCONNECTED_3831,
  SV2V_UNCONNECTED_3832,SV2V_UNCONNECTED_3833,SV2V_UNCONNECTED_3834,
  SV2V_UNCONNECTED_3835,SV2V_UNCONNECTED_3836,SV2V_UNCONNECTED_3837,
  SV2V_UNCONNECTED_3838,SV2V_UNCONNECTED_3839,SV2V_UNCONNECTED_3840,
  SV2V_UNCONNECTED_3841,SV2V_UNCONNECTED_3842,SV2V_UNCONNECTED_3843,
  SV2V_UNCONNECTED_3844,SV2V_UNCONNECTED_3845,SV2V_UNCONNECTED_3846,
  SV2V_UNCONNECTED_3847,SV2V_UNCONNECTED_3848,SV2V_UNCONNECTED_3849,
  SV2V_UNCONNECTED_3850,SV2V_UNCONNECTED_3851,SV2V_UNCONNECTED_3852,
  SV2V_UNCONNECTED_3853,SV2V_UNCONNECTED_3854,SV2V_UNCONNECTED_3855,
  SV2V_UNCONNECTED_3856,SV2V_UNCONNECTED_3857,SV2V_UNCONNECTED_3858,
  SV2V_UNCONNECTED_3859,SV2V_UNCONNECTED_3860,SV2V_UNCONNECTED_3861,
  SV2V_UNCONNECTED_3862,SV2V_UNCONNECTED_3863,SV2V_UNCONNECTED_3864,
  SV2V_UNCONNECTED_3865,SV2V_UNCONNECTED_3866,SV2V_UNCONNECTED_3867,SV2V_UNCONNECTED_3868,
  SV2V_UNCONNECTED_3869,SV2V_UNCONNECTED_3870,SV2V_UNCONNECTED_3871,
  SV2V_UNCONNECTED_3872,SV2V_UNCONNECTED_3873,SV2V_UNCONNECTED_3874,
  SV2V_UNCONNECTED_3875,SV2V_UNCONNECTED_3876,SV2V_UNCONNECTED_3877,
  SV2V_UNCONNECTED_3878,SV2V_UNCONNECTED_3879,SV2V_UNCONNECTED_3880,
  SV2V_UNCONNECTED_3881,SV2V_UNCONNECTED_3882,SV2V_UNCONNECTED_3883,
  SV2V_UNCONNECTED_3884,SV2V_UNCONNECTED_3885,SV2V_UNCONNECTED_3886,
  SV2V_UNCONNECTED_3887,SV2V_UNCONNECTED_3888,SV2V_UNCONNECTED_3889,
  SV2V_UNCONNECTED_3890,SV2V_UNCONNECTED_3891,SV2V_UNCONNECTED_3892,
  SV2V_UNCONNECTED_3893,SV2V_UNCONNECTED_3894,SV2V_UNCONNECTED_3895,
  SV2V_UNCONNECTED_3896,SV2V_UNCONNECTED_3897,SV2V_UNCONNECTED_3898,
  SV2V_UNCONNECTED_3899,SV2V_UNCONNECTED_3900,SV2V_UNCONNECTED_3901,
  SV2V_UNCONNECTED_3902,SV2V_UNCONNECTED_3903,SV2V_UNCONNECTED_3904,
  SV2V_UNCONNECTED_3905,SV2V_UNCONNECTED_3906,SV2V_UNCONNECTED_3907,SV2V_UNCONNECTED_3908,
  SV2V_UNCONNECTED_3909,SV2V_UNCONNECTED_3910,SV2V_UNCONNECTED_3911,
  SV2V_UNCONNECTED_3912,SV2V_UNCONNECTED_3913,SV2V_UNCONNECTED_3914,
  SV2V_UNCONNECTED_3915,SV2V_UNCONNECTED_3916,SV2V_UNCONNECTED_3917,
  SV2V_UNCONNECTED_3918,SV2V_UNCONNECTED_3919,SV2V_UNCONNECTED_3920,
  SV2V_UNCONNECTED_3921,SV2V_UNCONNECTED_3922,SV2V_UNCONNECTED_3923,
  SV2V_UNCONNECTED_3924,SV2V_UNCONNECTED_3925,SV2V_UNCONNECTED_3926,
  SV2V_UNCONNECTED_3927,SV2V_UNCONNECTED_3928,SV2V_UNCONNECTED_3929,
  SV2V_UNCONNECTED_3930,SV2V_UNCONNECTED_3931,SV2V_UNCONNECTED_3932,
  SV2V_UNCONNECTED_3933,SV2V_UNCONNECTED_3934,SV2V_UNCONNECTED_3935,
  SV2V_UNCONNECTED_3936,SV2V_UNCONNECTED_3937,SV2V_UNCONNECTED_3938,
  SV2V_UNCONNECTED_3939,SV2V_UNCONNECTED_3940,SV2V_UNCONNECTED_3941,
  SV2V_UNCONNECTED_3942,SV2V_UNCONNECTED_3943,SV2V_UNCONNECTED_3944,
  SV2V_UNCONNECTED_3945,SV2V_UNCONNECTED_3946,SV2V_UNCONNECTED_3947,SV2V_UNCONNECTED_3948,
  SV2V_UNCONNECTED_3949,SV2V_UNCONNECTED_3950,SV2V_UNCONNECTED_3951,
  SV2V_UNCONNECTED_3952,SV2V_UNCONNECTED_3953,SV2V_UNCONNECTED_3954,
  SV2V_UNCONNECTED_3955,SV2V_UNCONNECTED_3956,SV2V_UNCONNECTED_3957,
  SV2V_UNCONNECTED_3958,SV2V_UNCONNECTED_3959,SV2V_UNCONNECTED_3960,
  SV2V_UNCONNECTED_3961,SV2V_UNCONNECTED_3962,SV2V_UNCONNECTED_3963,
  SV2V_UNCONNECTED_3964,SV2V_UNCONNECTED_3965,SV2V_UNCONNECTED_3966,
  SV2V_UNCONNECTED_3967,SV2V_UNCONNECTED_3968,SV2V_UNCONNECTED_3969,
  SV2V_UNCONNECTED_3970,SV2V_UNCONNECTED_3971,SV2V_UNCONNECTED_3972,
  SV2V_UNCONNECTED_3973,SV2V_UNCONNECTED_3974,SV2V_UNCONNECTED_3975,
  SV2V_UNCONNECTED_3976,SV2V_UNCONNECTED_3977,SV2V_UNCONNECTED_3978,
  SV2V_UNCONNECTED_3979,SV2V_UNCONNECTED_3980,SV2V_UNCONNECTED_3981,
  SV2V_UNCONNECTED_3982,SV2V_UNCONNECTED_3983,SV2V_UNCONNECTED_3984,
  SV2V_UNCONNECTED_3985,SV2V_UNCONNECTED_3986,SV2V_UNCONNECTED_3987,SV2V_UNCONNECTED_3988,
  SV2V_UNCONNECTED_3989,SV2V_UNCONNECTED_3990,SV2V_UNCONNECTED_3991,
  SV2V_UNCONNECTED_3992,SV2V_UNCONNECTED_3993,SV2V_UNCONNECTED_3994,
  SV2V_UNCONNECTED_3995,SV2V_UNCONNECTED_3996,SV2V_UNCONNECTED_3997,
  SV2V_UNCONNECTED_3998,SV2V_UNCONNECTED_3999,SV2V_UNCONNECTED_4000,
  SV2V_UNCONNECTED_4001,SV2V_UNCONNECTED_4002,SV2V_UNCONNECTED_4003,
  SV2V_UNCONNECTED_4004,SV2V_UNCONNECTED_4005,SV2V_UNCONNECTED_4006,
  SV2V_UNCONNECTED_4007,SV2V_UNCONNECTED_4008,SV2V_UNCONNECTED_4009,
  SV2V_UNCONNECTED_4010,SV2V_UNCONNECTED_4011,SV2V_UNCONNECTED_4012,
  SV2V_UNCONNECTED_4013,SV2V_UNCONNECTED_4014,SV2V_UNCONNECTED_4015,
  SV2V_UNCONNECTED_4016,SV2V_UNCONNECTED_4017,SV2V_UNCONNECTED_4018,
  SV2V_UNCONNECTED_4019,SV2V_UNCONNECTED_4020,SV2V_UNCONNECTED_4021,
  SV2V_UNCONNECTED_4022,SV2V_UNCONNECTED_4023,SV2V_UNCONNECTED_4024,
  SV2V_UNCONNECTED_4025,SV2V_UNCONNECTED_4026,SV2V_UNCONNECTED_4027,SV2V_UNCONNECTED_4028,
  SV2V_UNCONNECTED_4029,SV2V_UNCONNECTED_4030,SV2V_UNCONNECTED_4031,
  SV2V_UNCONNECTED_4032,SV2V_UNCONNECTED_4033,SV2V_UNCONNECTED_4034,
  SV2V_UNCONNECTED_4035,SV2V_UNCONNECTED_4036,SV2V_UNCONNECTED_4037,
  SV2V_UNCONNECTED_4038,SV2V_UNCONNECTED_4039,SV2V_UNCONNECTED_4040,
  SV2V_UNCONNECTED_4041,SV2V_UNCONNECTED_4042,SV2V_UNCONNECTED_4043,
  SV2V_UNCONNECTED_4044,SV2V_UNCONNECTED_4045,SV2V_UNCONNECTED_4046,
  SV2V_UNCONNECTED_4047,SV2V_UNCONNECTED_4048,SV2V_UNCONNECTED_4049,
  SV2V_UNCONNECTED_4050,SV2V_UNCONNECTED_4051,SV2V_UNCONNECTED_4052,
  SV2V_UNCONNECTED_4053,SV2V_UNCONNECTED_4054,SV2V_UNCONNECTED_4055,
  SV2V_UNCONNECTED_4056,SV2V_UNCONNECTED_4057,SV2V_UNCONNECTED_4058,
  SV2V_UNCONNECTED_4059,SV2V_UNCONNECTED_4060,SV2V_UNCONNECTED_4061,
  SV2V_UNCONNECTED_4062,SV2V_UNCONNECTED_4063,SV2V_UNCONNECTED_4064,
  SV2V_UNCONNECTED_4065,SV2V_UNCONNECTED_4066,SV2V_UNCONNECTED_4067,SV2V_UNCONNECTED_4068,
  SV2V_UNCONNECTED_4069,SV2V_UNCONNECTED_4070,SV2V_UNCONNECTED_4071,
  SV2V_UNCONNECTED_4072,SV2V_UNCONNECTED_4073,SV2V_UNCONNECTED_4074,
  SV2V_UNCONNECTED_4075,SV2V_UNCONNECTED_4076,SV2V_UNCONNECTED_4077,
  SV2V_UNCONNECTED_4078,SV2V_UNCONNECTED_4079,SV2V_UNCONNECTED_4080,
  SV2V_UNCONNECTED_4081,SV2V_UNCONNECTED_4082,SV2V_UNCONNECTED_4083,
  SV2V_UNCONNECTED_4084,SV2V_UNCONNECTED_4085,SV2V_UNCONNECTED_4086,
  SV2V_UNCONNECTED_4087,SV2V_UNCONNECTED_4088,SV2V_UNCONNECTED_4089,
  SV2V_UNCONNECTED_4090,SV2V_UNCONNECTED_4091,SV2V_UNCONNECTED_4092,
  SV2V_UNCONNECTED_4093,SV2V_UNCONNECTED_4094,SV2V_UNCONNECTED_4095,
  SV2V_UNCONNECTED_4096,SV2V_UNCONNECTED_4097,SV2V_UNCONNECTED_4098,
  SV2V_UNCONNECTED_4099,SV2V_UNCONNECTED_4100,SV2V_UNCONNECTED_4101,
  SV2V_UNCONNECTED_4102,SV2V_UNCONNECTED_4103,SV2V_UNCONNECTED_4104,
  SV2V_UNCONNECTED_4105,SV2V_UNCONNECTED_4106,SV2V_UNCONNECTED_4107,SV2V_UNCONNECTED_4108,
  SV2V_UNCONNECTED_4109,SV2V_UNCONNECTED_4110,SV2V_UNCONNECTED_4111,
  SV2V_UNCONNECTED_4112,SV2V_UNCONNECTED_4113,SV2V_UNCONNECTED_4114,
  SV2V_UNCONNECTED_4115,SV2V_UNCONNECTED_4116,SV2V_UNCONNECTED_4117,
  SV2V_UNCONNECTED_4118,SV2V_UNCONNECTED_4119,SV2V_UNCONNECTED_4120,
  SV2V_UNCONNECTED_4121,SV2V_UNCONNECTED_4122,SV2V_UNCONNECTED_4123,
  SV2V_UNCONNECTED_4124,SV2V_UNCONNECTED_4125,SV2V_UNCONNECTED_4126,
  SV2V_UNCONNECTED_4127,SV2V_UNCONNECTED_4128,SV2V_UNCONNECTED_4129,
  SV2V_UNCONNECTED_4130,SV2V_UNCONNECTED_4131,SV2V_UNCONNECTED_4132,
  SV2V_UNCONNECTED_4133,SV2V_UNCONNECTED_4134,SV2V_UNCONNECTED_4135,
  SV2V_UNCONNECTED_4136,SV2V_UNCONNECTED_4137,SV2V_UNCONNECTED_4138,
  SV2V_UNCONNECTED_4139,SV2V_UNCONNECTED_4140,SV2V_UNCONNECTED_4141,
  SV2V_UNCONNECTED_4142,SV2V_UNCONNECTED_4143,SV2V_UNCONNECTED_4144,
  SV2V_UNCONNECTED_4145,SV2V_UNCONNECTED_4146,SV2V_UNCONNECTED_4147,SV2V_UNCONNECTED_4148,
  SV2V_UNCONNECTED_4149,SV2V_UNCONNECTED_4150,SV2V_UNCONNECTED_4151,
  SV2V_UNCONNECTED_4152,SV2V_UNCONNECTED_4153,SV2V_UNCONNECTED_4154,
  SV2V_UNCONNECTED_4155,SV2V_UNCONNECTED_4156,SV2V_UNCONNECTED_4157,
  SV2V_UNCONNECTED_4158,SV2V_UNCONNECTED_4159,SV2V_UNCONNECTED_4160,
  SV2V_UNCONNECTED_4161,SV2V_UNCONNECTED_4162,SV2V_UNCONNECTED_4163,
  SV2V_UNCONNECTED_4164,SV2V_UNCONNECTED_4165,SV2V_UNCONNECTED_4166,
  SV2V_UNCONNECTED_4167,SV2V_UNCONNECTED_4168,SV2V_UNCONNECTED_4169,
  SV2V_UNCONNECTED_4170,SV2V_UNCONNECTED_4171,SV2V_UNCONNECTED_4172,
  SV2V_UNCONNECTED_4173,SV2V_UNCONNECTED_4174,SV2V_UNCONNECTED_4175,
  SV2V_UNCONNECTED_4176,SV2V_UNCONNECTED_4177,SV2V_UNCONNECTED_4178,
  SV2V_UNCONNECTED_4179,SV2V_UNCONNECTED_4180,SV2V_UNCONNECTED_4181,
  SV2V_UNCONNECTED_4182,SV2V_UNCONNECTED_4183,SV2V_UNCONNECTED_4184,
  SV2V_UNCONNECTED_4185,SV2V_UNCONNECTED_4186,SV2V_UNCONNECTED_4187,SV2V_UNCONNECTED_4188,
  SV2V_UNCONNECTED_4189,SV2V_UNCONNECTED_4190,SV2V_UNCONNECTED_4191,
  SV2V_UNCONNECTED_4192,SV2V_UNCONNECTED_4193,SV2V_UNCONNECTED_4194,
  SV2V_UNCONNECTED_4195,SV2V_UNCONNECTED_4196,SV2V_UNCONNECTED_4197,
  SV2V_UNCONNECTED_4198,SV2V_UNCONNECTED_4199,SV2V_UNCONNECTED_4200,
  SV2V_UNCONNECTED_4201,SV2V_UNCONNECTED_4202,SV2V_UNCONNECTED_4203,
  SV2V_UNCONNECTED_4204,SV2V_UNCONNECTED_4205,SV2V_UNCONNECTED_4206,
  SV2V_UNCONNECTED_4207,SV2V_UNCONNECTED_4208,SV2V_UNCONNECTED_4209,
  SV2V_UNCONNECTED_4210,SV2V_UNCONNECTED_4211,SV2V_UNCONNECTED_4212,
  SV2V_UNCONNECTED_4213,SV2V_UNCONNECTED_4214,SV2V_UNCONNECTED_4215,
  SV2V_UNCONNECTED_4216,SV2V_UNCONNECTED_4217,SV2V_UNCONNECTED_4218,
  SV2V_UNCONNECTED_4219,SV2V_UNCONNECTED_4220,SV2V_UNCONNECTED_4221,
  SV2V_UNCONNECTED_4222,SV2V_UNCONNECTED_4223,SV2V_UNCONNECTED_4224,
  SV2V_UNCONNECTED_4225,SV2V_UNCONNECTED_4226,SV2V_UNCONNECTED_4227,SV2V_UNCONNECTED_4228,
  SV2V_UNCONNECTED_4229,SV2V_UNCONNECTED_4230,SV2V_UNCONNECTED_4231,
  SV2V_UNCONNECTED_4232,SV2V_UNCONNECTED_4233,SV2V_UNCONNECTED_4234,
  SV2V_UNCONNECTED_4235,SV2V_UNCONNECTED_4236,SV2V_UNCONNECTED_4237,
  SV2V_UNCONNECTED_4238,SV2V_UNCONNECTED_4239,SV2V_UNCONNECTED_4240,
  SV2V_UNCONNECTED_4241,SV2V_UNCONNECTED_4242,SV2V_UNCONNECTED_4243,
  SV2V_UNCONNECTED_4244,SV2V_UNCONNECTED_4245,SV2V_UNCONNECTED_4246,
  SV2V_UNCONNECTED_4247,SV2V_UNCONNECTED_4248,SV2V_UNCONNECTED_4249,
  SV2V_UNCONNECTED_4250,SV2V_UNCONNECTED_4251,SV2V_UNCONNECTED_4252,
  SV2V_UNCONNECTED_4253,SV2V_UNCONNECTED_4254,SV2V_UNCONNECTED_4255,
  SV2V_UNCONNECTED_4256,SV2V_UNCONNECTED_4257,SV2V_UNCONNECTED_4258,
  SV2V_UNCONNECTED_4259,SV2V_UNCONNECTED_4260,SV2V_UNCONNECTED_4261,
  SV2V_UNCONNECTED_4262,SV2V_UNCONNECTED_4263,SV2V_UNCONNECTED_4264,
  SV2V_UNCONNECTED_4265,SV2V_UNCONNECTED_4266,SV2V_UNCONNECTED_4267,SV2V_UNCONNECTED_4268,
  SV2V_UNCONNECTED_4269,SV2V_UNCONNECTED_4270,SV2V_UNCONNECTED_4271,
  SV2V_UNCONNECTED_4272,SV2V_UNCONNECTED_4273,SV2V_UNCONNECTED_4274,
  SV2V_UNCONNECTED_4275,SV2V_UNCONNECTED_4276,SV2V_UNCONNECTED_4277,
  SV2V_UNCONNECTED_4278,SV2V_UNCONNECTED_4279,SV2V_UNCONNECTED_4280,
  SV2V_UNCONNECTED_4281,SV2V_UNCONNECTED_4282,SV2V_UNCONNECTED_4283,
  SV2V_UNCONNECTED_4284,SV2V_UNCONNECTED_4285,SV2V_UNCONNECTED_4286,
  SV2V_UNCONNECTED_4287,SV2V_UNCONNECTED_4288,SV2V_UNCONNECTED_4289,
  SV2V_UNCONNECTED_4290,SV2V_UNCONNECTED_4291,SV2V_UNCONNECTED_4292,
  SV2V_UNCONNECTED_4293,SV2V_UNCONNECTED_4294,SV2V_UNCONNECTED_4295,
  SV2V_UNCONNECTED_4296,SV2V_UNCONNECTED_4297,SV2V_UNCONNECTED_4298,
  SV2V_UNCONNECTED_4299,SV2V_UNCONNECTED_4300,SV2V_UNCONNECTED_4301,
  SV2V_UNCONNECTED_4302,SV2V_UNCONNECTED_4303,SV2V_UNCONNECTED_4304,
  SV2V_UNCONNECTED_4305,SV2V_UNCONNECTED_4306,SV2V_UNCONNECTED_4307,SV2V_UNCONNECTED_4308,
  SV2V_UNCONNECTED_4309,SV2V_UNCONNECTED_4310,SV2V_UNCONNECTED_4311,
  SV2V_UNCONNECTED_4312,SV2V_UNCONNECTED_4313,SV2V_UNCONNECTED_4314,
  SV2V_UNCONNECTED_4315,SV2V_UNCONNECTED_4316,SV2V_UNCONNECTED_4317,
  SV2V_UNCONNECTED_4318,SV2V_UNCONNECTED_4319,SV2V_UNCONNECTED_4320,
  SV2V_UNCONNECTED_4321,SV2V_UNCONNECTED_4322,SV2V_UNCONNECTED_4323,
  SV2V_UNCONNECTED_4324,SV2V_UNCONNECTED_4325,SV2V_UNCONNECTED_4326,
  SV2V_UNCONNECTED_4327,SV2V_UNCONNECTED_4328,SV2V_UNCONNECTED_4329,
  SV2V_UNCONNECTED_4330,SV2V_UNCONNECTED_4331,SV2V_UNCONNECTED_4332,
  SV2V_UNCONNECTED_4333,SV2V_UNCONNECTED_4334,SV2V_UNCONNECTED_4335,
  SV2V_UNCONNECTED_4336,SV2V_UNCONNECTED_4337,SV2V_UNCONNECTED_4338,
  SV2V_UNCONNECTED_4339,SV2V_UNCONNECTED_4340,SV2V_UNCONNECTED_4341,
  SV2V_UNCONNECTED_4342,SV2V_UNCONNECTED_4343,SV2V_UNCONNECTED_4344,
  SV2V_UNCONNECTED_4345,SV2V_UNCONNECTED_4346,SV2V_UNCONNECTED_4347,SV2V_UNCONNECTED_4348,
  SV2V_UNCONNECTED_4349,SV2V_UNCONNECTED_4350,SV2V_UNCONNECTED_4351,
  SV2V_UNCONNECTED_4352,SV2V_UNCONNECTED_4353,SV2V_UNCONNECTED_4354,
  SV2V_UNCONNECTED_4355,SV2V_UNCONNECTED_4356,SV2V_UNCONNECTED_4357,
  SV2V_UNCONNECTED_4358,SV2V_UNCONNECTED_4359,SV2V_UNCONNECTED_4360,
  SV2V_UNCONNECTED_4361,SV2V_UNCONNECTED_4362,SV2V_UNCONNECTED_4363,
  SV2V_UNCONNECTED_4364,SV2V_UNCONNECTED_4365,SV2V_UNCONNECTED_4366,
  SV2V_UNCONNECTED_4367,SV2V_UNCONNECTED_4368,SV2V_UNCONNECTED_4369,
  SV2V_UNCONNECTED_4370,SV2V_UNCONNECTED_4371,SV2V_UNCONNECTED_4372,
  SV2V_UNCONNECTED_4373,SV2V_UNCONNECTED_4374,SV2V_UNCONNECTED_4375,
  SV2V_UNCONNECTED_4376,SV2V_UNCONNECTED_4377,SV2V_UNCONNECTED_4378,
  SV2V_UNCONNECTED_4379,SV2V_UNCONNECTED_4380,SV2V_UNCONNECTED_4381,
  SV2V_UNCONNECTED_4382,SV2V_UNCONNECTED_4383,SV2V_UNCONNECTED_4384,
  SV2V_UNCONNECTED_4385,SV2V_UNCONNECTED_4386,SV2V_UNCONNECTED_4387,SV2V_UNCONNECTED_4388,
  SV2V_UNCONNECTED_4389,SV2V_UNCONNECTED_4390,SV2V_UNCONNECTED_4391,
  SV2V_UNCONNECTED_4392,SV2V_UNCONNECTED_4393,SV2V_UNCONNECTED_4394,
  SV2V_UNCONNECTED_4395,SV2V_UNCONNECTED_4396,SV2V_UNCONNECTED_4397,
  SV2V_UNCONNECTED_4398,SV2V_UNCONNECTED_4399,SV2V_UNCONNECTED_4400,
  SV2V_UNCONNECTED_4401,SV2V_UNCONNECTED_4402,SV2V_UNCONNECTED_4403,
  SV2V_UNCONNECTED_4404,SV2V_UNCONNECTED_4405,SV2V_UNCONNECTED_4406,
  SV2V_UNCONNECTED_4407,SV2V_UNCONNECTED_4408,SV2V_UNCONNECTED_4409,
  SV2V_UNCONNECTED_4410,SV2V_UNCONNECTED_4411,SV2V_UNCONNECTED_4412,
  SV2V_UNCONNECTED_4413,SV2V_UNCONNECTED_4414,SV2V_UNCONNECTED_4415,
  SV2V_UNCONNECTED_4416,SV2V_UNCONNECTED_4417,SV2V_UNCONNECTED_4418,
  SV2V_UNCONNECTED_4419,SV2V_UNCONNECTED_4420,SV2V_UNCONNECTED_4421,
  SV2V_UNCONNECTED_4422,SV2V_UNCONNECTED_4423,SV2V_UNCONNECTED_4424,
  SV2V_UNCONNECTED_4425,SV2V_UNCONNECTED_4426,SV2V_UNCONNECTED_4427,SV2V_UNCONNECTED_4428,
  SV2V_UNCONNECTED_4429,SV2V_UNCONNECTED_4430,SV2V_UNCONNECTED_4431,
  SV2V_UNCONNECTED_4432,SV2V_UNCONNECTED_4433,SV2V_UNCONNECTED_4434,
  SV2V_UNCONNECTED_4435,SV2V_UNCONNECTED_4436,SV2V_UNCONNECTED_4437,
  SV2V_UNCONNECTED_4438,SV2V_UNCONNECTED_4439,SV2V_UNCONNECTED_4440,
  SV2V_UNCONNECTED_4441,SV2V_UNCONNECTED_4442,SV2V_UNCONNECTED_4443,
  SV2V_UNCONNECTED_4444,SV2V_UNCONNECTED_4445,SV2V_UNCONNECTED_4446,
  SV2V_UNCONNECTED_4447,SV2V_UNCONNECTED_4448,SV2V_UNCONNECTED_4449,
  SV2V_UNCONNECTED_4450,SV2V_UNCONNECTED_4451,SV2V_UNCONNECTED_4452,
  SV2V_UNCONNECTED_4453,SV2V_UNCONNECTED_4454,SV2V_UNCONNECTED_4455,
  SV2V_UNCONNECTED_4456,SV2V_UNCONNECTED_4457,SV2V_UNCONNECTED_4458,
  SV2V_UNCONNECTED_4459,SV2V_UNCONNECTED_4460,SV2V_UNCONNECTED_4461,
  SV2V_UNCONNECTED_4462,SV2V_UNCONNECTED_4463,SV2V_UNCONNECTED_4464,
  SV2V_UNCONNECTED_4465,SV2V_UNCONNECTED_4466,SV2V_UNCONNECTED_4467,SV2V_UNCONNECTED_4468,
  SV2V_UNCONNECTED_4469,SV2V_UNCONNECTED_4470,SV2V_UNCONNECTED_4471,
  SV2V_UNCONNECTED_4472,SV2V_UNCONNECTED_4473,SV2V_UNCONNECTED_4474,
  SV2V_UNCONNECTED_4475,SV2V_UNCONNECTED_4476,SV2V_UNCONNECTED_4477,
  SV2V_UNCONNECTED_4478,SV2V_UNCONNECTED_4479,SV2V_UNCONNECTED_4480,
  SV2V_UNCONNECTED_4481,SV2V_UNCONNECTED_4482,SV2V_UNCONNECTED_4483,
  SV2V_UNCONNECTED_4484,SV2V_UNCONNECTED_4485,SV2V_UNCONNECTED_4486,
  SV2V_UNCONNECTED_4487,SV2V_UNCONNECTED_4488,SV2V_UNCONNECTED_4489,
  SV2V_UNCONNECTED_4490,SV2V_UNCONNECTED_4491,SV2V_UNCONNECTED_4492,
  SV2V_UNCONNECTED_4493,SV2V_UNCONNECTED_4494,SV2V_UNCONNECTED_4495,
  SV2V_UNCONNECTED_4496,SV2V_UNCONNECTED_4497,SV2V_UNCONNECTED_4498,
  SV2V_UNCONNECTED_4499,SV2V_UNCONNECTED_4500,SV2V_UNCONNECTED_4501,
  SV2V_UNCONNECTED_4502,SV2V_UNCONNECTED_4503,SV2V_UNCONNECTED_4504,
  SV2V_UNCONNECTED_4505,SV2V_UNCONNECTED_4506,SV2V_UNCONNECTED_4507,SV2V_UNCONNECTED_4508,
  SV2V_UNCONNECTED_4509,SV2V_UNCONNECTED_4510,SV2V_UNCONNECTED_4511,
  SV2V_UNCONNECTED_4512,SV2V_UNCONNECTED_4513,SV2V_UNCONNECTED_4514,
  SV2V_UNCONNECTED_4515,SV2V_UNCONNECTED_4516,SV2V_UNCONNECTED_4517,
  SV2V_UNCONNECTED_4518,SV2V_UNCONNECTED_4519,SV2V_UNCONNECTED_4520,
  SV2V_UNCONNECTED_4521,SV2V_UNCONNECTED_4522,SV2V_UNCONNECTED_4523,
  SV2V_UNCONNECTED_4524,SV2V_UNCONNECTED_4525,SV2V_UNCONNECTED_4526,
  SV2V_UNCONNECTED_4527,SV2V_UNCONNECTED_4528,SV2V_UNCONNECTED_4529,
  SV2V_UNCONNECTED_4530,SV2V_UNCONNECTED_4531,SV2V_UNCONNECTED_4532,
  SV2V_UNCONNECTED_4533,SV2V_UNCONNECTED_4534,SV2V_UNCONNECTED_4535,
  SV2V_UNCONNECTED_4536,SV2V_UNCONNECTED_4537,SV2V_UNCONNECTED_4538,
  SV2V_UNCONNECTED_4539,SV2V_UNCONNECTED_4540,SV2V_UNCONNECTED_4541,
  SV2V_UNCONNECTED_4542,SV2V_UNCONNECTED_4543,SV2V_UNCONNECTED_4544,
  SV2V_UNCONNECTED_4545,SV2V_UNCONNECTED_4546,SV2V_UNCONNECTED_4547,SV2V_UNCONNECTED_4548,
  SV2V_UNCONNECTED_4549,SV2V_UNCONNECTED_4550,SV2V_UNCONNECTED_4551,
  SV2V_UNCONNECTED_4552,SV2V_UNCONNECTED_4553,SV2V_UNCONNECTED_4554,
  SV2V_UNCONNECTED_4555,SV2V_UNCONNECTED_4556,SV2V_UNCONNECTED_4557,
  SV2V_UNCONNECTED_4558,SV2V_UNCONNECTED_4559,SV2V_UNCONNECTED_4560,
  SV2V_UNCONNECTED_4561,SV2V_UNCONNECTED_4562,SV2V_UNCONNECTED_4563,
  SV2V_UNCONNECTED_4564,SV2V_UNCONNECTED_4565,SV2V_UNCONNECTED_4566,
  SV2V_UNCONNECTED_4567,SV2V_UNCONNECTED_4568,SV2V_UNCONNECTED_4569,
  SV2V_UNCONNECTED_4570,SV2V_UNCONNECTED_4571,SV2V_UNCONNECTED_4572,
  SV2V_UNCONNECTED_4573,SV2V_UNCONNECTED_4574,SV2V_UNCONNECTED_4575,
  SV2V_UNCONNECTED_4576,SV2V_UNCONNECTED_4577,SV2V_UNCONNECTED_4578,
  SV2V_UNCONNECTED_4579,SV2V_UNCONNECTED_4580,SV2V_UNCONNECTED_4581,
  SV2V_UNCONNECTED_4582,SV2V_UNCONNECTED_4583,SV2V_UNCONNECTED_4584,
  SV2V_UNCONNECTED_4585,SV2V_UNCONNECTED_4586,SV2V_UNCONNECTED_4587,SV2V_UNCONNECTED_4588,
  SV2V_UNCONNECTED_4589,SV2V_UNCONNECTED_4590,SV2V_UNCONNECTED_4591,
  SV2V_UNCONNECTED_4592,SV2V_UNCONNECTED_4593,SV2V_UNCONNECTED_4594,
  SV2V_UNCONNECTED_4595,SV2V_UNCONNECTED_4596,SV2V_UNCONNECTED_4597,
  SV2V_UNCONNECTED_4598,SV2V_UNCONNECTED_4599,SV2V_UNCONNECTED_4600,
  SV2V_UNCONNECTED_4601,SV2V_UNCONNECTED_4602,SV2V_UNCONNECTED_4603,
  SV2V_UNCONNECTED_4604,SV2V_UNCONNECTED_4605,SV2V_UNCONNECTED_4606,
  SV2V_UNCONNECTED_4607,SV2V_UNCONNECTED_4608,SV2V_UNCONNECTED_4609,
  SV2V_UNCONNECTED_4610,SV2V_UNCONNECTED_4611,SV2V_UNCONNECTED_4612,
  SV2V_UNCONNECTED_4613,SV2V_UNCONNECTED_4614,SV2V_UNCONNECTED_4615,
  SV2V_UNCONNECTED_4616,SV2V_UNCONNECTED_4617,SV2V_UNCONNECTED_4618,
  SV2V_UNCONNECTED_4619,SV2V_UNCONNECTED_4620,SV2V_UNCONNECTED_4621,
  SV2V_UNCONNECTED_4622,SV2V_UNCONNECTED_4623,SV2V_UNCONNECTED_4624,
  SV2V_UNCONNECTED_4625,SV2V_UNCONNECTED_4626,SV2V_UNCONNECTED_4627,SV2V_UNCONNECTED_4628,
  SV2V_UNCONNECTED_4629,SV2V_UNCONNECTED_4630,SV2V_UNCONNECTED_4631,
  SV2V_UNCONNECTED_4632,SV2V_UNCONNECTED_4633,SV2V_UNCONNECTED_4634,
  SV2V_UNCONNECTED_4635,SV2V_UNCONNECTED_4636,SV2V_UNCONNECTED_4637,
  SV2V_UNCONNECTED_4638,SV2V_UNCONNECTED_4639,SV2V_UNCONNECTED_4640,
  SV2V_UNCONNECTED_4641,SV2V_UNCONNECTED_4642,SV2V_UNCONNECTED_4643,
  SV2V_UNCONNECTED_4644,SV2V_UNCONNECTED_4645,SV2V_UNCONNECTED_4646,
  SV2V_UNCONNECTED_4647,SV2V_UNCONNECTED_4648,SV2V_UNCONNECTED_4649,
  SV2V_UNCONNECTED_4650,SV2V_UNCONNECTED_4651,SV2V_UNCONNECTED_4652,
  SV2V_UNCONNECTED_4653,SV2V_UNCONNECTED_4654,SV2V_UNCONNECTED_4655,
  SV2V_UNCONNECTED_4656,SV2V_UNCONNECTED_4657,SV2V_UNCONNECTED_4658,
  SV2V_UNCONNECTED_4659,SV2V_UNCONNECTED_4660,SV2V_UNCONNECTED_4661,
  SV2V_UNCONNECTED_4662,SV2V_UNCONNECTED_4663,SV2V_UNCONNECTED_4664,
  SV2V_UNCONNECTED_4665,SV2V_UNCONNECTED_4666,SV2V_UNCONNECTED_4667,SV2V_UNCONNECTED_4668,
  SV2V_UNCONNECTED_4669,SV2V_UNCONNECTED_4670,SV2V_UNCONNECTED_4671,
  SV2V_UNCONNECTED_4672,SV2V_UNCONNECTED_4673,SV2V_UNCONNECTED_4674,
  SV2V_UNCONNECTED_4675,SV2V_UNCONNECTED_4676,SV2V_UNCONNECTED_4677,
  SV2V_UNCONNECTED_4678,SV2V_UNCONNECTED_4679,SV2V_UNCONNECTED_4680,
  SV2V_UNCONNECTED_4681,SV2V_UNCONNECTED_4682,SV2V_UNCONNECTED_4683,
  SV2V_UNCONNECTED_4684,SV2V_UNCONNECTED_4685,SV2V_UNCONNECTED_4686,
  SV2V_UNCONNECTED_4687,SV2V_UNCONNECTED_4688,SV2V_UNCONNECTED_4689,
  SV2V_UNCONNECTED_4690,SV2V_UNCONNECTED_4691,SV2V_UNCONNECTED_4692,
  SV2V_UNCONNECTED_4693,SV2V_UNCONNECTED_4694,SV2V_UNCONNECTED_4695,
  SV2V_UNCONNECTED_4696,SV2V_UNCONNECTED_4697,SV2V_UNCONNECTED_4698,
  SV2V_UNCONNECTED_4699,SV2V_UNCONNECTED_4700,SV2V_UNCONNECTED_4701,
  SV2V_UNCONNECTED_4702,SV2V_UNCONNECTED_4703,SV2V_UNCONNECTED_4704,
  SV2V_UNCONNECTED_4705,SV2V_UNCONNECTED_4706,SV2V_UNCONNECTED_4707,SV2V_UNCONNECTED_4708,
  SV2V_UNCONNECTED_4709,SV2V_UNCONNECTED_4710,SV2V_UNCONNECTED_4711,
  SV2V_UNCONNECTED_4712,SV2V_UNCONNECTED_4713,SV2V_UNCONNECTED_4714,
  SV2V_UNCONNECTED_4715,SV2V_UNCONNECTED_4716,SV2V_UNCONNECTED_4717,
  SV2V_UNCONNECTED_4718,SV2V_UNCONNECTED_4719,SV2V_UNCONNECTED_4720,
  SV2V_UNCONNECTED_4721,SV2V_UNCONNECTED_4722,SV2V_UNCONNECTED_4723,
  SV2V_UNCONNECTED_4724,SV2V_UNCONNECTED_4725,SV2V_UNCONNECTED_4726,
  SV2V_UNCONNECTED_4727,SV2V_UNCONNECTED_4728,SV2V_UNCONNECTED_4729,
  SV2V_UNCONNECTED_4730,SV2V_UNCONNECTED_4731,SV2V_UNCONNECTED_4732,
  SV2V_UNCONNECTED_4733,SV2V_UNCONNECTED_4734,SV2V_UNCONNECTED_4735,
  SV2V_UNCONNECTED_4736,SV2V_UNCONNECTED_4737,SV2V_UNCONNECTED_4738,
  SV2V_UNCONNECTED_4739,SV2V_UNCONNECTED_4740,SV2V_UNCONNECTED_4741,
  SV2V_UNCONNECTED_4742,SV2V_UNCONNECTED_4743,SV2V_UNCONNECTED_4744,
  SV2V_UNCONNECTED_4745,SV2V_UNCONNECTED_4746,SV2V_UNCONNECTED_4747,SV2V_UNCONNECTED_4748,
  SV2V_UNCONNECTED_4749,SV2V_UNCONNECTED_4750,SV2V_UNCONNECTED_4751,
  SV2V_UNCONNECTED_4752,SV2V_UNCONNECTED_4753,SV2V_UNCONNECTED_4754,
  SV2V_UNCONNECTED_4755,SV2V_UNCONNECTED_4756,SV2V_UNCONNECTED_4757,
  SV2V_UNCONNECTED_4758,SV2V_UNCONNECTED_4759,SV2V_UNCONNECTED_4760,
  SV2V_UNCONNECTED_4761,SV2V_UNCONNECTED_4762,SV2V_UNCONNECTED_4763,
  SV2V_UNCONNECTED_4764,SV2V_UNCONNECTED_4765,SV2V_UNCONNECTED_4766,
  SV2V_UNCONNECTED_4767,SV2V_UNCONNECTED_4768,SV2V_UNCONNECTED_4769,
  SV2V_UNCONNECTED_4770,SV2V_UNCONNECTED_4771,SV2V_UNCONNECTED_4772,
  SV2V_UNCONNECTED_4773,SV2V_UNCONNECTED_4774,SV2V_UNCONNECTED_4775,
  SV2V_UNCONNECTED_4776,SV2V_UNCONNECTED_4777,SV2V_UNCONNECTED_4778,
  SV2V_UNCONNECTED_4779,SV2V_UNCONNECTED_4780,SV2V_UNCONNECTED_4781,
  SV2V_UNCONNECTED_4782,SV2V_UNCONNECTED_4783,SV2V_UNCONNECTED_4784,
  SV2V_UNCONNECTED_4785,SV2V_UNCONNECTED_4786,SV2V_UNCONNECTED_4787,SV2V_UNCONNECTED_4788,
  SV2V_UNCONNECTED_4789,SV2V_UNCONNECTED_4790,SV2V_UNCONNECTED_4791,
  SV2V_UNCONNECTED_4792,SV2V_UNCONNECTED_4793,SV2V_UNCONNECTED_4794,
  SV2V_UNCONNECTED_4795,SV2V_UNCONNECTED_4796,SV2V_UNCONNECTED_4797,
  SV2V_UNCONNECTED_4798,SV2V_UNCONNECTED_4799,SV2V_UNCONNECTED_4800,
  SV2V_UNCONNECTED_4801,SV2V_UNCONNECTED_4802,SV2V_UNCONNECTED_4803,
  SV2V_UNCONNECTED_4804,SV2V_UNCONNECTED_4805,SV2V_UNCONNECTED_4806,
  SV2V_UNCONNECTED_4807,SV2V_UNCONNECTED_4808,SV2V_UNCONNECTED_4809,
  SV2V_UNCONNECTED_4810,SV2V_UNCONNECTED_4811,SV2V_UNCONNECTED_4812,
  SV2V_UNCONNECTED_4813,SV2V_UNCONNECTED_4814,SV2V_UNCONNECTED_4815,
  SV2V_UNCONNECTED_4816,SV2V_UNCONNECTED_4817,SV2V_UNCONNECTED_4818,
  SV2V_UNCONNECTED_4819,SV2V_UNCONNECTED_4820,SV2V_UNCONNECTED_4821,
  SV2V_UNCONNECTED_4822,SV2V_UNCONNECTED_4823,SV2V_UNCONNECTED_4824,
  SV2V_UNCONNECTED_4825,SV2V_UNCONNECTED_4826,SV2V_UNCONNECTED_4827,SV2V_UNCONNECTED_4828,
  SV2V_UNCONNECTED_4829,SV2V_UNCONNECTED_4830,SV2V_UNCONNECTED_4831,
  SV2V_UNCONNECTED_4832,SV2V_UNCONNECTED_4833,SV2V_UNCONNECTED_4834,
  SV2V_UNCONNECTED_4835,SV2V_UNCONNECTED_4836,SV2V_UNCONNECTED_4837,
  SV2V_UNCONNECTED_4838,SV2V_UNCONNECTED_4839,SV2V_UNCONNECTED_4840,
  SV2V_UNCONNECTED_4841,SV2V_UNCONNECTED_4842,SV2V_UNCONNECTED_4843,
  SV2V_UNCONNECTED_4844,SV2V_UNCONNECTED_4845,SV2V_UNCONNECTED_4846,
  SV2V_UNCONNECTED_4847,SV2V_UNCONNECTED_4848,SV2V_UNCONNECTED_4849,
  SV2V_UNCONNECTED_4850,SV2V_UNCONNECTED_4851,SV2V_UNCONNECTED_4852,
  SV2V_UNCONNECTED_4853,SV2V_UNCONNECTED_4854,SV2V_UNCONNECTED_4855,
  SV2V_UNCONNECTED_4856,SV2V_UNCONNECTED_4857,SV2V_UNCONNECTED_4858,
  SV2V_UNCONNECTED_4859,SV2V_UNCONNECTED_4860,SV2V_UNCONNECTED_4861,
  SV2V_UNCONNECTED_4862,SV2V_UNCONNECTED_4863,SV2V_UNCONNECTED_4864,
  SV2V_UNCONNECTED_4865,SV2V_UNCONNECTED_4866,SV2V_UNCONNECTED_4867,SV2V_UNCONNECTED_4868,
  SV2V_UNCONNECTED_4869,SV2V_UNCONNECTED_4870,SV2V_UNCONNECTED_4871,
  SV2V_UNCONNECTED_4872,SV2V_UNCONNECTED_4873,SV2V_UNCONNECTED_4874,
  SV2V_UNCONNECTED_4875,SV2V_UNCONNECTED_4876,SV2V_UNCONNECTED_4877,
  SV2V_UNCONNECTED_4878,SV2V_UNCONNECTED_4879,SV2V_UNCONNECTED_4880,
  SV2V_UNCONNECTED_4881,SV2V_UNCONNECTED_4882,SV2V_UNCONNECTED_4883,
  SV2V_UNCONNECTED_4884,SV2V_UNCONNECTED_4885,SV2V_UNCONNECTED_4886,
  SV2V_UNCONNECTED_4887,SV2V_UNCONNECTED_4888,SV2V_UNCONNECTED_4889,
  SV2V_UNCONNECTED_4890,SV2V_UNCONNECTED_4891,SV2V_UNCONNECTED_4892,
  SV2V_UNCONNECTED_4893,SV2V_UNCONNECTED_4894,SV2V_UNCONNECTED_4895,
  SV2V_UNCONNECTED_4896,SV2V_UNCONNECTED_4897,SV2V_UNCONNECTED_4898,
  SV2V_UNCONNECTED_4899,SV2V_UNCONNECTED_4900,SV2V_UNCONNECTED_4901,
  SV2V_UNCONNECTED_4902,SV2V_UNCONNECTED_4903,SV2V_UNCONNECTED_4904,
  SV2V_UNCONNECTED_4905,SV2V_UNCONNECTED_4906,SV2V_UNCONNECTED_4907,SV2V_UNCONNECTED_4908,
  SV2V_UNCONNECTED_4909,SV2V_UNCONNECTED_4910,SV2V_UNCONNECTED_4911,
  SV2V_UNCONNECTED_4912,SV2V_UNCONNECTED_4913,SV2V_UNCONNECTED_4914,
  SV2V_UNCONNECTED_4915,SV2V_UNCONNECTED_4916,SV2V_UNCONNECTED_4917,
  SV2V_UNCONNECTED_4918,SV2V_UNCONNECTED_4919,SV2V_UNCONNECTED_4920,
  SV2V_UNCONNECTED_4921,SV2V_UNCONNECTED_4922,SV2V_UNCONNECTED_4923,
  SV2V_UNCONNECTED_4924,SV2V_UNCONNECTED_4925,SV2V_UNCONNECTED_4926,
  SV2V_UNCONNECTED_4927,SV2V_UNCONNECTED_4928,SV2V_UNCONNECTED_4929,
  SV2V_UNCONNECTED_4930,SV2V_UNCONNECTED_4931,SV2V_UNCONNECTED_4932,
  SV2V_UNCONNECTED_4933,SV2V_UNCONNECTED_4934,SV2V_UNCONNECTED_4935,
  SV2V_UNCONNECTED_4936,SV2V_UNCONNECTED_4937,SV2V_UNCONNECTED_4938,
  SV2V_UNCONNECTED_4939,SV2V_UNCONNECTED_4940,SV2V_UNCONNECTED_4941,
  SV2V_UNCONNECTED_4942,SV2V_UNCONNECTED_4943,SV2V_UNCONNECTED_4944,
  SV2V_UNCONNECTED_4945,SV2V_UNCONNECTED_4946,SV2V_UNCONNECTED_4947,SV2V_UNCONNECTED_4948,
  SV2V_UNCONNECTED_4949,SV2V_UNCONNECTED_4950,SV2V_UNCONNECTED_4951,
  SV2V_UNCONNECTED_4952,SV2V_UNCONNECTED_4953,SV2V_UNCONNECTED_4954,
  SV2V_UNCONNECTED_4955,SV2V_UNCONNECTED_4956,SV2V_UNCONNECTED_4957,
  SV2V_UNCONNECTED_4958,SV2V_UNCONNECTED_4959,SV2V_UNCONNECTED_4960,
  SV2V_UNCONNECTED_4961,SV2V_UNCONNECTED_4962,SV2V_UNCONNECTED_4963,
  SV2V_UNCONNECTED_4964,SV2V_UNCONNECTED_4965,SV2V_UNCONNECTED_4966,
  SV2V_UNCONNECTED_4967,SV2V_UNCONNECTED_4968,SV2V_UNCONNECTED_4969,
  SV2V_UNCONNECTED_4970,SV2V_UNCONNECTED_4971,SV2V_UNCONNECTED_4972,
  SV2V_UNCONNECTED_4973,SV2V_UNCONNECTED_4974,SV2V_UNCONNECTED_4975,
  SV2V_UNCONNECTED_4976,SV2V_UNCONNECTED_4977,SV2V_UNCONNECTED_4978,
  SV2V_UNCONNECTED_4979,SV2V_UNCONNECTED_4980,SV2V_UNCONNECTED_4981,
  SV2V_UNCONNECTED_4982,SV2V_UNCONNECTED_4983,SV2V_UNCONNECTED_4984,
  SV2V_UNCONNECTED_4985,SV2V_UNCONNECTED_4986,SV2V_UNCONNECTED_4987,SV2V_UNCONNECTED_4988,
  SV2V_UNCONNECTED_4989,SV2V_UNCONNECTED_4990,SV2V_UNCONNECTED_4991,
  SV2V_UNCONNECTED_4992,SV2V_UNCONNECTED_4993,SV2V_UNCONNECTED_4994,
  SV2V_UNCONNECTED_4995,SV2V_UNCONNECTED_4996,SV2V_UNCONNECTED_4997,
  SV2V_UNCONNECTED_4998,SV2V_UNCONNECTED_4999,SV2V_UNCONNECTED_5000,
  SV2V_UNCONNECTED_5001,SV2V_UNCONNECTED_5002,SV2V_UNCONNECTED_5003,
  SV2V_UNCONNECTED_5004,SV2V_UNCONNECTED_5005,SV2V_UNCONNECTED_5006,
  SV2V_UNCONNECTED_5007,SV2V_UNCONNECTED_5008,SV2V_UNCONNECTED_5009,
  SV2V_UNCONNECTED_5010,SV2V_UNCONNECTED_5011,SV2V_UNCONNECTED_5012,
  SV2V_UNCONNECTED_5013,SV2V_UNCONNECTED_5014,SV2V_UNCONNECTED_5015,
  SV2V_UNCONNECTED_5016,SV2V_UNCONNECTED_5017,SV2V_UNCONNECTED_5018,
  SV2V_UNCONNECTED_5019,SV2V_UNCONNECTED_5020,SV2V_UNCONNECTED_5021,
  SV2V_UNCONNECTED_5022,SV2V_UNCONNECTED_5023,SV2V_UNCONNECTED_5024,
  SV2V_UNCONNECTED_5025,SV2V_UNCONNECTED_5026,SV2V_UNCONNECTED_5027,SV2V_UNCONNECTED_5028,
  SV2V_UNCONNECTED_5029,SV2V_UNCONNECTED_5030,SV2V_UNCONNECTED_5031,
  SV2V_UNCONNECTED_5032,SV2V_UNCONNECTED_5033,SV2V_UNCONNECTED_5034,
  SV2V_UNCONNECTED_5035,SV2V_UNCONNECTED_5036,SV2V_UNCONNECTED_5037,
  SV2V_UNCONNECTED_5038,SV2V_UNCONNECTED_5039,SV2V_UNCONNECTED_5040,
  SV2V_UNCONNECTED_5041,SV2V_UNCONNECTED_5042,SV2V_UNCONNECTED_5043,
  SV2V_UNCONNECTED_5044,SV2V_UNCONNECTED_5045,SV2V_UNCONNECTED_5046,
  SV2V_UNCONNECTED_5047,SV2V_UNCONNECTED_5048,SV2V_UNCONNECTED_5049,
  SV2V_UNCONNECTED_5050,SV2V_UNCONNECTED_5051,SV2V_UNCONNECTED_5052,
  SV2V_UNCONNECTED_5053,SV2V_UNCONNECTED_5054,SV2V_UNCONNECTED_5055,
  SV2V_UNCONNECTED_5056,SV2V_UNCONNECTED_5057,SV2V_UNCONNECTED_5058,
  SV2V_UNCONNECTED_5059,SV2V_UNCONNECTED_5060,SV2V_UNCONNECTED_5061,
  SV2V_UNCONNECTED_5062,SV2V_UNCONNECTED_5063,SV2V_UNCONNECTED_5064,
  SV2V_UNCONNECTED_5065,SV2V_UNCONNECTED_5066,SV2V_UNCONNECTED_5067,SV2V_UNCONNECTED_5068,
  SV2V_UNCONNECTED_5069,SV2V_UNCONNECTED_5070,SV2V_UNCONNECTED_5071,
  SV2V_UNCONNECTED_5072,SV2V_UNCONNECTED_5073,SV2V_UNCONNECTED_5074,
  SV2V_UNCONNECTED_5075,SV2V_UNCONNECTED_5076,SV2V_UNCONNECTED_5077,
  SV2V_UNCONNECTED_5078,SV2V_UNCONNECTED_5079,SV2V_UNCONNECTED_5080,
  SV2V_UNCONNECTED_5081,SV2V_UNCONNECTED_5082,SV2V_UNCONNECTED_5083,
  SV2V_UNCONNECTED_5084,SV2V_UNCONNECTED_5085,SV2V_UNCONNECTED_5086,
  SV2V_UNCONNECTED_5087,SV2V_UNCONNECTED_5088,SV2V_UNCONNECTED_5089,
  SV2V_UNCONNECTED_5090,SV2V_UNCONNECTED_5091,SV2V_UNCONNECTED_5092,
  SV2V_UNCONNECTED_5093,SV2V_UNCONNECTED_5094,SV2V_UNCONNECTED_5095,
  SV2V_UNCONNECTED_5096,SV2V_UNCONNECTED_5097,SV2V_UNCONNECTED_5098,
  SV2V_UNCONNECTED_5099,SV2V_UNCONNECTED_5100,SV2V_UNCONNECTED_5101,
  SV2V_UNCONNECTED_5102,SV2V_UNCONNECTED_5103,SV2V_UNCONNECTED_5104,
  SV2V_UNCONNECTED_5105,SV2V_UNCONNECTED_5106,SV2V_UNCONNECTED_5107,SV2V_UNCONNECTED_5108,
  SV2V_UNCONNECTED_5109,SV2V_UNCONNECTED_5110,SV2V_UNCONNECTED_5111,
  SV2V_UNCONNECTED_5112,SV2V_UNCONNECTED_5113,SV2V_UNCONNECTED_5114,
  SV2V_UNCONNECTED_5115,SV2V_UNCONNECTED_5116,SV2V_UNCONNECTED_5117,
  SV2V_UNCONNECTED_5118,SV2V_UNCONNECTED_5119,SV2V_UNCONNECTED_5120,
  SV2V_UNCONNECTED_5121,SV2V_UNCONNECTED_5122,SV2V_UNCONNECTED_5123,
  SV2V_UNCONNECTED_5124,SV2V_UNCONNECTED_5125,SV2V_UNCONNECTED_5126,
  SV2V_UNCONNECTED_5127,SV2V_UNCONNECTED_5128,SV2V_UNCONNECTED_5129,
  SV2V_UNCONNECTED_5130,SV2V_UNCONNECTED_5131,SV2V_UNCONNECTED_5132,
  SV2V_UNCONNECTED_5133,SV2V_UNCONNECTED_5134,SV2V_UNCONNECTED_5135,
  SV2V_UNCONNECTED_5136,SV2V_UNCONNECTED_5137,SV2V_UNCONNECTED_5138,
  SV2V_UNCONNECTED_5139,SV2V_UNCONNECTED_5140,SV2V_UNCONNECTED_5141,
  SV2V_UNCONNECTED_5142,SV2V_UNCONNECTED_5143,SV2V_UNCONNECTED_5144,
  SV2V_UNCONNECTED_5145,SV2V_UNCONNECTED_5146,SV2V_UNCONNECTED_5147,SV2V_UNCONNECTED_5148,
  SV2V_UNCONNECTED_5149,SV2V_UNCONNECTED_5150,SV2V_UNCONNECTED_5151,
  SV2V_UNCONNECTED_5152,SV2V_UNCONNECTED_5153,SV2V_UNCONNECTED_5154,
  SV2V_UNCONNECTED_5155,SV2V_UNCONNECTED_5156,SV2V_UNCONNECTED_5157,
  SV2V_UNCONNECTED_5158,SV2V_UNCONNECTED_5159,SV2V_UNCONNECTED_5160,
  SV2V_UNCONNECTED_5161,SV2V_UNCONNECTED_5162,SV2V_UNCONNECTED_5163,
  SV2V_UNCONNECTED_5164,SV2V_UNCONNECTED_5165,SV2V_UNCONNECTED_5166,
  SV2V_UNCONNECTED_5167,SV2V_UNCONNECTED_5168,SV2V_UNCONNECTED_5169,
  SV2V_UNCONNECTED_5170,SV2V_UNCONNECTED_5171,SV2V_UNCONNECTED_5172,
  SV2V_UNCONNECTED_5173,SV2V_UNCONNECTED_5174,SV2V_UNCONNECTED_5175,
  SV2V_UNCONNECTED_5176,SV2V_UNCONNECTED_5177,SV2V_UNCONNECTED_5178,
  SV2V_UNCONNECTED_5179,SV2V_UNCONNECTED_5180,SV2V_UNCONNECTED_5181,
  SV2V_UNCONNECTED_5182,SV2V_UNCONNECTED_5183,SV2V_UNCONNECTED_5184,
  SV2V_UNCONNECTED_5185,SV2V_UNCONNECTED_5186,SV2V_UNCONNECTED_5187,SV2V_UNCONNECTED_5188,
  SV2V_UNCONNECTED_5189,SV2V_UNCONNECTED_5190,SV2V_UNCONNECTED_5191,
  SV2V_UNCONNECTED_5192,SV2V_UNCONNECTED_5193,SV2V_UNCONNECTED_5194,
  SV2V_UNCONNECTED_5195,SV2V_UNCONNECTED_5196,SV2V_UNCONNECTED_5197,
  SV2V_UNCONNECTED_5198,SV2V_UNCONNECTED_5199,SV2V_UNCONNECTED_5200,
  SV2V_UNCONNECTED_5201,SV2V_UNCONNECTED_5202,SV2V_UNCONNECTED_5203,
  SV2V_UNCONNECTED_5204,SV2V_UNCONNECTED_5205,SV2V_UNCONNECTED_5206,
  SV2V_UNCONNECTED_5207,SV2V_UNCONNECTED_5208,SV2V_UNCONNECTED_5209,
  SV2V_UNCONNECTED_5210,SV2V_UNCONNECTED_5211,SV2V_UNCONNECTED_5212,
  SV2V_UNCONNECTED_5213,SV2V_UNCONNECTED_5214,SV2V_UNCONNECTED_5215,
  SV2V_UNCONNECTED_5216,SV2V_UNCONNECTED_5217,SV2V_UNCONNECTED_5218,
  SV2V_UNCONNECTED_5219,SV2V_UNCONNECTED_5220,SV2V_UNCONNECTED_5221,
  SV2V_UNCONNECTED_5222,SV2V_UNCONNECTED_5223,SV2V_UNCONNECTED_5224,
  SV2V_UNCONNECTED_5225,SV2V_UNCONNECTED_5226,SV2V_UNCONNECTED_5227,SV2V_UNCONNECTED_5228,
  SV2V_UNCONNECTED_5229,SV2V_UNCONNECTED_5230,SV2V_UNCONNECTED_5231,
  SV2V_UNCONNECTED_5232,SV2V_UNCONNECTED_5233,SV2V_UNCONNECTED_5234,
  SV2V_UNCONNECTED_5235,SV2V_UNCONNECTED_5236,SV2V_UNCONNECTED_5237,
  SV2V_UNCONNECTED_5238,SV2V_UNCONNECTED_5239,SV2V_UNCONNECTED_5240,
  SV2V_UNCONNECTED_5241,SV2V_UNCONNECTED_5242,SV2V_UNCONNECTED_5243,
  SV2V_UNCONNECTED_5244,SV2V_UNCONNECTED_5245,SV2V_UNCONNECTED_5246,
  SV2V_UNCONNECTED_5247,SV2V_UNCONNECTED_5248,SV2V_UNCONNECTED_5249,
  SV2V_UNCONNECTED_5250,SV2V_UNCONNECTED_5251,SV2V_UNCONNECTED_5252,
  SV2V_UNCONNECTED_5253,SV2V_UNCONNECTED_5254,SV2V_UNCONNECTED_5255,
  SV2V_UNCONNECTED_5256,SV2V_UNCONNECTED_5257,SV2V_UNCONNECTED_5258,
  SV2V_UNCONNECTED_5259,SV2V_UNCONNECTED_5260,SV2V_UNCONNECTED_5261,
  SV2V_UNCONNECTED_5262,SV2V_UNCONNECTED_5263,SV2V_UNCONNECTED_5264,
  SV2V_UNCONNECTED_5265,SV2V_UNCONNECTED_5266,SV2V_UNCONNECTED_5267,SV2V_UNCONNECTED_5268,
  SV2V_UNCONNECTED_5269,SV2V_UNCONNECTED_5270,SV2V_UNCONNECTED_5271,
  SV2V_UNCONNECTED_5272,SV2V_UNCONNECTED_5273,SV2V_UNCONNECTED_5274,
  SV2V_UNCONNECTED_5275,SV2V_UNCONNECTED_5276,SV2V_UNCONNECTED_5277,
  SV2V_UNCONNECTED_5278,SV2V_UNCONNECTED_5279,SV2V_UNCONNECTED_5280,
  SV2V_UNCONNECTED_5281,SV2V_UNCONNECTED_5282,SV2V_UNCONNECTED_5283,
  SV2V_UNCONNECTED_5284,SV2V_UNCONNECTED_5285,SV2V_UNCONNECTED_5286,
  SV2V_UNCONNECTED_5287,SV2V_UNCONNECTED_5288,SV2V_UNCONNECTED_5289,
  SV2V_UNCONNECTED_5290,SV2V_UNCONNECTED_5291,SV2V_UNCONNECTED_5292,
  SV2V_UNCONNECTED_5293,SV2V_UNCONNECTED_5294,SV2V_UNCONNECTED_5295,
  SV2V_UNCONNECTED_5296,SV2V_UNCONNECTED_5297,SV2V_UNCONNECTED_5298,
  SV2V_UNCONNECTED_5299,SV2V_UNCONNECTED_5300,SV2V_UNCONNECTED_5301,
  SV2V_UNCONNECTED_5302,SV2V_UNCONNECTED_5303,SV2V_UNCONNECTED_5304,
  SV2V_UNCONNECTED_5305,SV2V_UNCONNECTED_5306,SV2V_UNCONNECTED_5307,SV2V_UNCONNECTED_5308,
  SV2V_UNCONNECTED_5309,SV2V_UNCONNECTED_5310,SV2V_UNCONNECTED_5311,
  SV2V_UNCONNECTED_5312,SV2V_UNCONNECTED_5313,SV2V_UNCONNECTED_5314,
  SV2V_UNCONNECTED_5315,SV2V_UNCONNECTED_5316,SV2V_UNCONNECTED_5317,
  SV2V_UNCONNECTED_5318,SV2V_UNCONNECTED_5319,SV2V_UNCONNECTED_5320,
  SV2V_UNCONNECTED_5321,SV2V_UNCONNECTED_5322,SV2V_UNCONNECTED_5323,
  SV2V_UNCONNECTED_5324,SV2V_UNCONNECTED_5325,SV2V_UNCONNECTED_5326,
  SV2V_UNCONNECTED_5327,SV2V_UNCONNECTED_5328,SV2V_UNCONNECTED_5329,
  SV2V_UNCONNECTED_5330,SV2V_UNCONNECTED_5331,SV2V_UNCONNECTED_5332,
  SV2V_UNCONNECTED_5333,SV2V_UNCONNECTED_5334,SV2V_UNCONNECTED_5335,
  SV2V_UNCONNECTED_5336,SV2V_UNCONNECTED_5337,SV2V_UNCONNECTED_5338,
  SV2V_UNCONNECTED_5339,SV2V_UNCONNECTED_5340,SV2V_UNCONNECTED_5341,
  SV2V_UNCONNECTED_5342,SV2V_UNCONNECTED_5343,SV2V_UNCONNECTED_5344,
  SV2V_UNCONNECTED_5345,SV2V_UNCONNECTED_5346,SV2V_UNCONNECTED_5347,SV2V_UNCONNECTED_5348,
  SV2V_UNCONNECTED_5349,SV2V_UNCONNECTED_5350,SV2V_UNCONNECTED_5351,
  SV2V_UNCONNECTED_5352,SV2V_UNCONNECTED_5353,SV2V_UNCONNECTED_5354,
  SV2V_UNCONNECTED_5355,SV2V_UNCONNECTED_5356,SV2V_UNCONNECTED_5357,
  SV2V_UNCONNECTED_5358,SV2V_UNCONNECTED_5359,SV2V_UNCONNECTED_5360,
  SV2V_UNCONNECTED_5361,SV2V_UNCONNECTED_5362,SV2V_UNCONNECTED_5363,
  SV2V_UNCONNECTED_5364,SV2V_UNCONNECTED_5365,SV2V_UNCONNECTED_5366,
  SV2V_UNCONNECTED_5367,SV2V_UNCONNECTED_5368,SV2V_UNCONNECTED_5369,
  SV2V_UNCONNECTED_5370,SV2V_UNCONNECTED_5371,SV2V_UNCONNECTED_5372,
  SV2V_UNCONNECTED_5373,SV2V_UNCONNECTED_5374,SV2V_UNCONNECTED_5375,
  SV2V_UNCONNECTED_5376,SV2V_UNCONNECTED_5377,SV2V_UNCONNECTED_5378,
  SV2V_UNCONNECTED_5379,SV2V_UNCONNECTED_5380,SV2V_UNCONNECTED_5381,
  SV2V_UNCONNECTED_5382,SV2V_UNCONNECTED_5383,SV2V_UNCONNECTED_5384,
  SV2V_UNCONNECTED_5385,SV2V_UNCONNECTED_5386,SV2V_UNCONNECTED_5387,SV2V_UNCONNECTED_5388,
  SV2V_UNCONNECTED_5389,SV2V_UNCONNECTED_5390,SV2V_UNCONNECTED_5391,
  SV2V_UNCONNECTED_5392,SV2V_UNCONNECTED_5393,SV2V_UNCONNECTED_5394,
  SV2V_UNCONNECTED_5395,SV2V_UNCONNECTED_5396,SV2V_UNCONNECTED_5397,
  SV2V_UNCONNECTED_5398,SV2V_UNCONNECTED_5399,SV2V_UNCONNECTED_5400,
  SV2V_UNCONNECTED_5401,SV2V_UNCONNECTED_5402,SV2V_UNCONNECTED_5403,
  SV2V_UNCONNECTED_5404,SV2V_UNCONNECTED_5405,SV2V_UNCONNECTED_5406,
  SV2V_UNCONNECTED_5407,SV2V_UNCONNECTED_5408,SV2V_UNCONNECTED_5409,
  SV2V_UNCONNECTED_5410,SV2V_UNCONNECTED_5411,SV2V_UNCONNECTED_5412,
  SV2V_UNCONNECTED_5413,SV2V_UNCONNECTED_5414,SV2V_UNCONNECTED_5415,
  SV2V_UNCONNECTED_5416,SV2V_UNCONNECTED_5417,SV2V_UNCONNECTED_5418,
  SV2V_UNCONNECTED_5419,SV2V_UNCONNECTED_5420,SV2V_UNCONNECTED_5421,
  SV2V_UNCONNECTED_5422,SV2V_UNCONNECTED_5423,SV2V_UNCONNECTED_5424,
  SV2V_UNCONNECTED_5425,SV2V_UNCONNECTED_5426,SV2V_UNCONNECTED_5427,SV2V_UNCONNECTED_5428,
  SV2V_UNCONNECTED_5429,SV2V_UNCONNECTED_5430,SV2V_UNCONNECTED_5431,
  SV2V_UNCONNECTED_5432,SV2V_UNCONNECTED_5433,SV2V_UNCONNECTED_5434,
  SV2V_UNCONNECTED_5435,SV2V_UNCONNECTED_5436,SV2V_UNCONNECTED_5437,
  SV2V_UNCONNECTED_5438,SV2V_UNCONNECTED_5439,SV2V_UNCONNECTED_5440,
  SV2V_UNCONNECTED_5441,SV2V_UNCONNECTED_5442,SV2V_UNCONNECTED_5443,
  SV2V_UNCONNECTED_5444,SV2V_UNCONNECTED_5445,SV2V_UNCONNECTED_5446,
  SV2V_UNCONNECTED_5447,SV2V_UNCONNECTED_5448,SV2V_UNCONNECTED_5449,
  SV2V_UNCONNECTED_5450,SV2V_UNCONNECTED_5451,SV2V_UNCONNECTED_5452,
  SV2V_UNCONNECTED_5453,SV2V_UNCONNECTED_5454,SV2V_UNCONNECTED_5455,
  SV2V_UNCONNECTED_5456,SV2V_UNCONNECTED_5457,SV2V_UNCONNECTED_5458,
  SV2V_UNCONNECTED_5459,SV2V_UNCONNECTED_5460,SV2V_UNCONNECTED_5461,
  SV2V_UNCONNECTED_5462,SV2V_UNCONNECTED_5463,SV2V_UNCONNECTED_5464,
  SV2V_UNCONNECTED_5465,SV2V_UNCONNECTED_5466,SV2V_UNCONNECTED_5467,SV2V_UNCONNECTED_5468,
  SV2V_UNCONNECTED_5469,SV2V_UNCONNECTED_5470,SV2V_UNCONNECTED_5471,
  SV2V_UNCONNECTED_5472,SV2V_UNCONNECTED_5473,SV2V_UNCONNECTED_5474,
  SV2V_UNCONNECTED_5475,SV2V_UNCONNECTED_5476,SV2V_UNCONNECTED_5477,
  SV2V_UNCONNECTED_5478,SV2V_UNCONNECTED_5479,SV2V_UNCONNECTED_5480,
  SV2V_UNCONNECTED_5481,SV2V_UNCONNECTED_5482,SV2V_UNCONNECTED_5483,
  SV2V_UNCONNECTED_5484,SV2V_UNCONNECTED_5485,SV2V_UNCONNECTED_5486,
  SV2V_UNCONNECTED_5487,SV2V_UNCONNECTED_5488,SV2V_UNCONNECTED_5489,
  SV2V_UNCONNECTED_5490,SV2V_UNCONNECTED_5491,SV2V_UNCONNECTED_5492,
  SV2V_UNCONNECTED_5493,SV2V_UNCONNECTED_5494,SV2V_UNCONNECTED_5495,
  SV2V_UNCONNECTED_5496,SV2V_UNCONNECTED_5497,SV2V_UNCONNECTED_5498,
  SV2V_UNCONNECTED_5499,SV2V_UNCONNECTED_5500,SV2V_UNCONNECTED_5501,
  SV2V_UNCONNECTED_5502,SV2V_UNCONNECTED_5503,SV2V_UNCONNECTED_5504,
  SV2V_UNCONNECTED_5505,SV2V_UNCONNECTED_5506,SV2V_UNCONNECTED_5507,SV2V_UNCONNECTED_5508,
  SV2V_UNCONNECTED_5509,SV2V_UNCONNECTED_5510,SV2V_UNCONNECTED_5511,
  SV2V_UNCONNECTED_5512,SV2V_UNCONNECTED_5513,SV2V_UNCONNECTED_5514,
  SV2V_UNCONNECTED_5515,SV2V_UNCONNECTED_5516,SV2V_UNCONNECTED_5517,
  SV2V_UNCONNECTED_5518,SV2V_UNCONNECTED_5519,SV2V_UNCONNECTED_5520,
  SV2V_UNCONNECTED_5521,SV2V_UNCONNECTED_5522,SV2V_UNCONNECTED_5523,
  SV2V_UNCONNECTED_5524,SV2V_UNCONNECTED_5525,SV2V_UNCONNECTED_5526,
  SV2V_UNCONNECTED_5527,SV2V_UNCONNECTED_5528,SV2V_UNCONNECTED_5529,
  SV2V_UNCONNECTED_5530,SV2V_UNCONNECTED_5531,SV2V_UNCONNECTED_5532,
  SV2V_UNCONNECTED_5533,SV2V_UNCONNECTED_5534,SV2V_UNCONNECTED_5535,
  SV2V_UNCONNECTED_5536,SV2V_UNCONNECTED_5537,SV2V_UNCONNECTED_5538,
  SV2V_UNCONNECTED_5539,SV2V_UNCONNECTED_5540,SV2V_UNCONNECTED_5541,
  SV2V_UNCONNECTED_5542,SV2V_UNCONNECTED_5543,SV2V_UNCONNECTED_5544,
  SV2V_UNCONNECTED_5545,SV2V_UNCONNECTED_5546,SV2V_UNCONNECTED_5547,SV2V_UNCONNECTED_5548,
  SV2V_UNCONNECTED_5549,SV2V_UNCONNECTED_5550,SV2V_UNCONNECTED_5551,
  SV2V_UNCONNECTED_5552,SV2V_UNCONNECTED_5553,SV2V_UNCONNECTED_5554,
  SV2V_UNCONNECTED_5555,SV2V_UNCONNECTED_5556,SV2V_UNCONNECTED_5557,
  SV2V_UNCONNECTED_5558,SV2V_UNCONNECTED_5559,SV2V_UNCONNECTED_5560,
  SV2V_UNCONNECTED_5561,SV2V_UNCONNECTED_5562,SV2V_UNCONNECTED_5563,
  SV2V_UNCONNECTED_5564,SV2V_UNCONNECTED_5565,SV2V_UNCONNECTED_5566,
  SV2V_UNCONNECTED_5567,SV2V_UNCONNECTED_5568,SV2V_UNCONNECTED_5569,
  SV2V_UNCONNECTED_5570,SV2V_UNCONNECTED_5571,SV2V_UNCONNECTED_5572,
  SV2V_UNCONNECTED_5573,SV2V_UNCONNECTED_5574,SV2V_UNCONNECTED_5575,
  SV2V_UNCONNECTED_5576,SV2V_UNCONNECTED_5577,SV2V_UNCONNECTED_5578,
  SV2V_UNCONNECTED_5579,SV2V_UNCONNECTED_5580,SV2V_UNCONNECTED_5581,
  SV2V_UNCONNECTED_5582,SV2V_UNCONNECTED_5583,SV2V_UNCONNECTED_5584,
  SV2V_UNCONNECTED_5585,SV2V_UNCONNECTED_5586,SV2V_UNCONNECTED_5587,SV2V_UNCONNECTED_5588,
  SV2V_UNCONNECTED_5589,SV2V_UNCONNECTED_5590,SV2V_UNCONNECTED_5591,
  SV2V_UNCONNECTED_5592,SV2V_UNCONNECTED_5593,SV2V_UNCONNECTED_5594,
  SV2V_UNCONNECTED_5595,SV2V_UNCONNECTED_5596,SV2V_UNCONNECTED_5597,
  SV2V_UNCONNECTED_5598,SV2V_UNCONNECTED_5599,SV2V_UNCONNECTED_5600,
  SV2V_UNCONNECTED_5601,SV2V_UNCONNECTED_5602,SV2V_UNCONNECTED_5603,
  SV2V_UNCONNECTED_5604,SV2V_UNCONNECTED_5605,SV2V_UNCONNECTED_5606,
  SV2V_UNCONNECTED_5607,SV2V_UNCONNECTED_5608,SV2V_UNCONNECTED_5609,
  SV2V_UNCONNECTED_5610,SV2V_UNCONNECTED_5611,SV2V_UNCONNECTED_5612,
  SV2V_UNCONNECTED_5613,SV2V_UNCONNECTED_5614,SV2V_UNCONNECTED_5615,
  SV2V_UNCONNECTED_5616,SV2V_UNCONNECTED_5617,SV2V_UNCONNECTED_5618,
  SV2V_UNCONNECTED_5619,SV2V_UNCONNECTED_5620,SV2V_UNCONNECTED_5621,
  SV2V_UNCONNECTED_5622,SV2V_UNCONNECTED_5623,SV2V_UNCONNECTED_5624,
  SV2V_UNCONNECTED_5625,SV2V_UNCONNECTED_5626,SV2V_UNCONNECTED_5627,SV2V_UNCONNECTED_5628,
  SV2V_UNCONNECTED_5629,SV2V_UNCONNECTED_5630,SV2V_UNCONNECTED_5631,
  SV2V_UNCONNECTED_5632,SV2V_UNCONNECTED_5633,SV2V_UNCONNECTED_5634,
  SV2V_UNCONNECTED_5635,SV2V_UNCONNECTED_5636,SV2V_UNCONNECTED_5637,
  SV2V_UNCONNECTED_5638,SV2V_UNCONNECTED_5639,SV2V_UNCONNECTED_5640,
  SV2V_UNCONNECTED_5641,SV2V_UNCONNECTED_5642,SV2V_UNCONNECTED_5643,
  SV2V_UNCONNECTED_5644,SV2V_UNCONNECTED_5645,SV2V_UNCONNECTED_5646,
  SV2V_UNCONNECTED_5647,SV2V_UNCONNECTED_5648,SV2V_UNCONNECTED_5649,
  SV2V_UNCONNECTED_5650,SV2V_UNCONNECTED_5651,SV2V_UNCONNECTED_5652,
  SV2V_UNCONNECTED_5653,SV2V_UNCONNECTED_5654,SV2V_UNCONNECTED_5655,
  SV2V_UNCONNECTED_5656,SV2V_UNCONNECTED_5657,SV2V_UNCONNECTED_5658,
  SV2V_UNCONNECTED_5659,SV2V_UNCONNECTED_5660,SV2V_UNCONNECTED_5661,
  SV2V_UNCONNECTED_5662,SV2V_UNCONNECTED_5663,SV2V_UNCONNECTED_5664,
  SV2V_UNCONNECTED_5665,SV2V_UNCONNECTED_5666,SV2V_UNCONNECTED_5667,SV2V_UNCONNECTED_5668,
  SV2V_UNCONNECTED_5669,SV2V_UNCONNECTED_5670,SV2V_UNCONNECTED_5671,
  SV2V_UNCONNECTED_5672,SV2V_UNCONNECTED_5673,SV2V_UNCONNECTED_5674,
  SV2V_UNCONNECTED_5675,SV2V_UNCONNECTED_5676,SV2V_UNCONNECTED_5677,
  SV2V_UNCONNECTED_5678,SV2V_UNCONNECTED_5679,SV2V_UNCONNECTED_5680,
  SV2V_UNCONNECTED_5681,SV2V_UNCONNECTED_5682,SV2V_UNCONNECTED_5683,
  SV2V_UNCONNECTED_5684,SV2V_UNCONNECTED_5685,SV2V_UNCONNECTED_5686,
  SV2V_UNCONNECTED_5687,SV2V_UNCONNECTED_5688,SV2V_UNCONNECTED_5689,
  SV2V_UNCONNECTED_5690,SV2V_UNCONNECTED_5691,SV2V_UNCONNECTED_5692,
  SV2V_UNCONNECTED_5693,SV2V_UNCONNECTED_5694,SV2V_UNCONNECTED_5695,
  SV2V_UNCONNECTED_5696,SV2V_UNCONNECTED_5697,SV2V_UNCONNECTED_5698,
  SV2V_UNCONNECTED_5699,SV2V_UNCONNECTED_5700,SV2V_UNCONNECTED_5701,
  SV2V_UNCONNECTED_5702,SV2V_UNCONNECTED_5703,SV2V_UNCONNECTED_5704,
  SV2V_UNCONNECTED_5705,SV2V_UNCONNECTED_5706,SV2V_UNCONNECTED_5707,SV2V_UNCONNECTED_5708,
  SV2V_UNCONNECTED_5709,SV2V_UNCONNECTED_5710,SV2V_UNCONNECTED_5711,
  SV2V_UNCONNECTED_5712,SV2V_UNCONNECTED_5713,SV2V_UNCONNECTED_5714,
  SV2V_UNCONNECTED_5715,SV2V_UNCONNECTED_5716,SV2V_UNCONNECTED_5717,
  SV2V_UNCONNECTED_5718,SV2V_UNCONNECTED_5719,SV2V_UNCONNECTED_5720,
  SV2V_UNCONNECTED_5721,SV2V_UNCONNECTED_5722,SV2V_UNCONNECTED_5723,
  SV2V_UNCONNECTED_5724,SV2V_UNCONNECTED_5725,SV2V_UNCONNECTED_5726,
  SV2V_UNCONNECTED_5727,SV2V_UNCONNECTED_5728,SV2V_UNCONNECTED_5729,
  SV2V_UNCONNECTED_5730,SV2V_UNCONNECTED_5731,SV2V_UNCONNECTED_5732,
  SV2V_UNCONNECTED_5733,SV2V_UNCONNECTED_5734,SV2V_UNCONNECTED_5735,
  SV2V_UNCONNECTED_5736,SV2V_UNCONNECTED_5737,SV2V_UNCONNECTED_5738,
  SV2V_UNCONNECTED_5739,SV2V_UNCONNECTED_5740,SV2V_UNCONNECTED_5741,
  SV2V_UNCONNECTED_5742,SV2V_UNCONNECTED_5743,SV2V_UNCONNECTED_5744,
  SV2V_UNCONNECTED_5745,SV2V_UNCONNECTED_5746,SV2V_UNCONNECTED_5747,SV2V_UNCONNECTED_5748,
  SV2V_UNCONNECTED_5749,SV2V_UNCONNECTED_5750,SV2V_UNCONNECTED_5751,
  SV2V_UNCONNECTED_5752,SV2V_UNCONNECTED_5753,SV2V_UNCONNECTED_5754,
  SV2V_UNCONNECTED_5755,SV2V_UNCONNECTED_5756,SV2V_UNCONNECTED_5757,
  SV2V_UNCONNECTED_5758,SV2V_UNCONNECTED_5759,SV2V_UNCONNECTED_5760,
  SV2V_UNCONNECTED_5761,SV2V_UNCONNECTED_5762,SV2V_UNCONNECTED_5763,
  SV2V_UNCONNECTED_5764,SV2V_UNCONNECTED_5765,SV2V_UNCONNECTED_5766,
  SV2V_UNCONNECTED_5767,SV2V_UNCONNECTED_5768,SV2V_UNCONNECTED_5769,
  SV2V_UNCONNECTED_5770,SV2V_UNCONNECTED_5771,SV2V_UNCONNECTED_5772,
  SV2V_UNCONNECTED_5773,SV2V_UNCONNECTED_5774,SV2V_UNCONNECTED_5775,
  SV2V_UNCONNECTED_5776,SV2V_UNCONNECTED_5777,SV2V_UNCONNECTED_5778,
  SV2V_UNCONNECTED_5779,SV2V_UNCONNECTED_5780,SV2V_UNCONNECTED_5781,
  SV2V_UNCONNECTED_5782,SV2V_UNCONNECTED_5783,SV2V_UNCONNECTED_5784,
  SV2V_UNCONNECTED_5785,SV2V_UNCONNECTED_5786,SV2V_UNCONNECTED_5787,SV2V_UNCONNECTED_5788,
  SV2V_UNCONNECTED_5789,SV2V_UNCONNECTED_5790,SV2V_UNCONNECTED_5791,
  SV2V_UNCONNECTED_5792,SV2V_UNCONNECTED_5793,SV2V_UNCONNECTED_5794,
  SV2V_UNCONNECTED_5795,SV2V_UNCONNECTED_5796,SV2V_UNCONNECTED_5797,
  SV2V_UNCONNECTED_5798,SV2V_UNCONNECTED_5799,SV2V_UNCONNECTED_5800,
  SV2V_UNCONNECTED_5801,SV2V_UNCONNECTED_5802,SV2V_UNCONNECTED_5803,
  SV2V_UNCONNECTED_5804,SV2V_UNCONNECTED_5805,SV2V_UNCONNECTED_5806,
  SV2V_UNCONNECTED_5807,SV2V_UNCONNECTED_5808,SV2V_UNCONNECTED_5809,
  SV2V_UNCONNECTED_5810,SV2V_UNCONNECTED_5811,SV2V_UNCONNECTED_5812,
  SV2V_UNCONNECTED_5813,SV2V_UNCONNECTED_5814,SV2V_UNCONNECTED_5815,
  SV2V_UNCONNECTED_5816,SV2V_UNCONNECTED_5817,SV2V_UNCONNECTED_5818,
  SV2V_UNCONNECTED_5819,SV2V_UNCONNECTED_5820,SV2V_UNCONNECTED_5821,
  SV2V_UNCONNECTED_5822,SV2V_UNCONNECTED_5823,SV2V_UNCONNECTED_5824,
  SV2V_UNCONNECTED_5825,SV2V_UNCONNECTED_5826,SV2V_UNCONNECTED_5827,SV2V_UNCONNECTED_5828,
  SV2V_UNCONNECTED_5829,SV2V_UNCONNECTED_5830,SV2V_UNCONNECTED_5831,
  SV2V_UNCONNECTED_5832,SV2V_UNCONNECTED_5833,SV2V_UNCONNECTED_5834,
  SV2V_UNCONNECTED_5835,SV2V_UNCONNECTED_5836,SV2V_UNCONNECTED_5837,
  SV2V_UNCONNECTED_5838,SV2V_UNCONNECTED_5839,SV2V_UNCONNECTED_5840,
  SV2V_UNCONNECTED_5841,SV2V_UNCONNECTED_5842,SV2V_UNCONNECTED_5843,
  SV2V_UNCONNECTED_5844,SV2V_UNCONNECTED_5845,SV2V_UNCONNECTED_5846,
  SV2V_UNCONNECTED_5847,SV2V_UNCONNECTED_5848,SV2V_UNCONNECTED_5849,
  SV2V_UNCONNECTED_5850,SV2V_UNCONNECTED_5851,SV2V_UNCONNECTED_5852,
  SV2V_UNCONNECTED_5853,SV2V_UNCONNECTED_5854,SV2V_UNCONNECTED_5855,
  SV2V_UNCONNECTED_5856,SV2V_UNCONNECTED_5857,SV2V_UNCONNECTED_5858,
  SV2V_UNCONNECTED_5859,SV2V_UNCONNECTED_5860,SV2V_UNCONNECTED_5861,
  SV2V_UNCONNECTED_5862,SV2V_UNCONNECTED_5863,SV2V_UNCONNECTED_5864,
  SV2V_UNCONNECTED_5865,SV2V_UNCONNECTED_5866,SV2V_UNCONNECTED_5867,SV2V_UNCONNECTED_5868,
  SV2V_UNCONNECTED_5869,SV2V_UNCONNECTED_5870,SV2V_UNCONNECTED_5871,
  SV2V_UNCONNECTED_5872,SV2V_UNCONNECTED_5873,SV2V_UNCONNECTED_5874,
  SV2V_UNCONNECTED_5875,SV2V_UNCONNECTED_5876,SV2V_UNCONNECTED_5877,
  SV2V_UNCONNECTED_5878,SV2V_UNCONNECTED_5879,SV2V_UNCONNECTED_5880,
  SV2V_UNCONNECTED_5881,SV2V_UNCONNECTED_5882,SV2V_UNCONNECTED_5883,
  SV2V_UNCONNECTED_5884,SV2V_UNCONNECTED_5885,SV2V_UNCONNECTED_5886,
  SV2V_UNCONNECTED_5887,SV2V_UNCONNECTED_5888,SV2V_UNCONNECTED_5889,
  SV2V_UNCONNECTED_5890,SV2V_UNCONNECTED_5891,SV2V_UNCONNECTED_5892,
  SV2V_UNCONNECTED_5893,SV2V_UNCONNECTED_5894,SV2V_UNCONNECTED_5895,
  SV2V_UNCONNECTED_5896,SV2V_UNCONNECTED_5897,SV2V_UNCONNECTED_5898,
  SV2V_UNCONNECTED_5899,SV2V_UNCONNECTED_5900,SV2V_UNCONNECTED_5901,
  SV2V_UNCONNECTED_5902,SV2V_UNCONNECTED_5903,SV2V_UNCONNECTED_5904,
  SV2V_UNCONNECTED_5905,SV2V_UNCONNECTED_5906,SV2V_UNCONNECTED_5907,SV2V_UNCONNECTED_5908,
  SV2V_UNCONNECTED_5909,SV2V_UNCONNECTED_5910,SV2V_UNCONNECTED_5911,
  SV2V_UNCONNECTED_5912,SV2V_UNCONNECTED_5913,SV2V_UNCONNECTED_5914,
  SV2V_UNCONNECTED_5915,SV2V_UNCONNECTED_5916,SV2V_UNCONNECTED_5917,
  SV2V_UNCONNECTED_5918,SV2V_UNCONNECTED_5919,SV2V_UNCONNECTED_5920,
  SV2V_UNCONNECTED_5921,SV2V_UNCONNECTED_5922,SV2V_UNCONNECTED_5923,
  SV2V_UNCONNECTED_5924,SV2V_UNCONNECTED_5925,SV2V_UNCONNECTED_5926,
  SV2V_UNCONNECTED_5927,SV2V_UNCONNECTED_5928,SV2V_UNCONNECTED_5929,
  SV2V_UNCONNECTED_5930,SV2V_UNCONNECTED_5931,SV2V_UNCONNECTED_5932,
  SV2V_UNCONNECTED_5933,SV2V_UNCONNECTED_5934,SV2V_UNCONNECTED_5935,
  SV2V_UNCONNECTED_5936,SV2V_UNCONNECTED_5937,SV2V_UNCONNECTED_5938,
  SV2V_UNCONNECTED_5939,SV2V_UNCONNECTED_5940,SV2V_UNCONNECTED_5941,
  SV2V_UNCONNECTED_5942,SV2V_UNCONNECTED_5943,SV2V_UNCONNECTED_5944,
  SV2V_UNCONNECTED_5945,SV2V_UNCONNECTED_5946,SV2V_UNCONNECTED_5947,SV2V_UNCONNECTED_5948,
  SV2V_UNCONNECTED_5949,SV2V_UNCONNECTED_5950,SV2V_UNCONNECTED_5951,
  SV2V_UNCONNECTED_5952,SV2V_UNCONNECTED_5953,SV2V_UNCONNECTED_5954,
  SV2V_UNCONNECTED_5955,SV2V_UNCONNECTED_5956,SV2V_UNCONNECTED_5957,
  SV2V_UNCONNECTED_5958,SV2V_UNCONNECTED_5959,SV2V_UNCONNECTED_5960,
  SV2V_UNCONNECTED_5961,SV2V_UNCONNECTED_5962,SV2V_UNCONNECTED_5963,
  SV2V_UNCONNECTED_5964,SV2V_UNCONNECTED_5965,SV2V_UNCONNECTED_5966,
  SV2V_UNCONNECTED_5967,SV2V_UNCONNECTED_5968,SV2V_UNCONNECTED_5969,
  SV2V_UNCONNECTED_5970,SV2V_UNCONNECTED_5971,SV2V_UNCONNECTED_5972,
  SV2V_UNCONNECTED_5973,SV2V_UNCONNECTED_5974,SV2V_UNCONNECTED_5975,
  SV2V_UNCONNECTED_5976,SV2V_UNCONNECTED_5977,SV2V_UNCONNECTED_5978,
  SV2V_UNCONNECTED_5979,SV2V_UNCONNECTED_5980,SV2V_UNCONNECTED_5981,
  SV2V_UNCONNECTED_5982,SV2V_UNCONNECTED_5983,SV2V_UNCONNECTED_5984,
  SV2V_UNCONNECTED_5985,SV2V_UNCONNECTED_5986,SV2V_UNCONNECTED_5987,SV2V_UNCONNECTED_5988,
  SV2V_UNCONNECTED_5989,SV2V_UNCONNECTED_5990,SV2V_UNCONNECTED_5991,
  SV2V_UNCONNECTED_5992,SV2V_UNCONNECTED_5993,SV2V_UNCONNECTED_5994,
  SV2V_UNCONNECTED_5995,SV2V_UNCONNECTED_5996,SV2V_UNCONNECTED_5997,
  SV2V_UNCONNECTED_5998,SV2V_UNCONNECTED_5999,SV2V_UNCONNECTED_6000,
  SV2V_UNCONNECTED_6001,SV2V_UNCONNECTED_6002,SV2V_UNCONNECTED_6003,
  SV2V_UNCONNECTED_6004,SV2V_UNCONNECTED_6005,SV2V_UNCONNECTED_6006,
  SV2V_UNCONNECTED_6007,SV2V_UNCONNECTED_6008,SV2V_UNCONNECTED_6009,
  SV2V_UNCONNECTED_6010,SV2V_UNCONNECTED_6011,SV2V_UNCONNECTED_6012,
  SV2V_UNCONNECTED_6013,SV2V_UNCONNECTED_6014,SV2V_UNCONNECTED_6015,
  SV2V_UNCONNECTED_6016,SV2V_UNCONNECTED_6017,SV2V_UNCONNECTED_6018,
  SV2V_UNCONNECTED_6019,SV2V_UNCONNECTED_6020,SV2V_UNCONNECTED_6021,
  SV2V_UNCONNECTED_6022,SV2V_UNCONNECTED_6023,SV2V_UNCONNECTED_6024,
  SV2V_UNCONNECTED_6025,SV2V_UNCONNECTED_6026,SV2V_UNCONNECTED_6027,SV2V_UNCONNECTED_6028,
  SV2V_UNCONNECTED_6029,SV2V_UNCONNECTED_6030,SV2V_UNCONNECTED_6031,
  SV2V_UNCONNECTED_6032,SV2V_UNCONNECTED_6033,SV2V_UNCONNECTED_6034,
  SV2V_UNCONNECTED_6035,SV2V_UNCONNECTED_6036,SV2V_UNCONNECTED_6037,
  SV2V_UNCONNECTED_6038,SV2V_UNCONNECTED_6039,SV2V_UNCONNECTED_6040,
  SV2V_UNCONNECTED_6041,SV2V_UNCONNECTED_6042,SV2V_UNCONNECTED_6043,
  SV2V_UNCONNECTED_6044,SV2V_UNCONNECTED_6045,SV2V_UNCONNECTED_6046,
  SV2V_UNCONNECTED_6047,SV2V_UNCONNECTED_6048,SV2V_UNCONNECTED_6049,
  SV2V_UNCONNECTED_6050,SV2V_UNCONNECTED_6051,SV2V_UNCONNECTED_6052,
  SV2V_UNCONNECTED_6053,SV2V_UNCONNECTED_6054,SV2V_UNCONNECTED_6055,
  SV2V_UNCONNECTED_6056,SV2V_UNCONNECTED_6057,SV2V_UNCONNECTED_6058,
  SV2V_UNCONNECTED_6059,SV2V_UNCONNECTED_6060,SV2V_UNCONNECTED_6061,
  SV2V_UNCONNECTED_6062,SV2V_UNCONNECTED_6063,SV2V_UNCONNECTED_6064,
  SV2V_UNCONNECTED_6065,SV2V_UNCONNECTED_6066,SV2V_UNCONNECTED_6067,SV2V_UNCONNECTED_6068,
  SV2V_UNCONNECTED_6069,SV2V_UNCONNECTED_6070,SV2V_UNCONNECTED_6071,
  SV2V_UNCONNECTED_6072,SV2V_UNCONNECTED_6073,SV2V_UNCONNECTED_6074,
  SV2V_UNCONNECTED_6075,SV2V_UNCONNECTED_6076,SV2V_UNCONNECTED_6077,
  SV2V_UNCONNECTED_6078,SV2V_UNCONNECTED_6079,SV2V_UNCONNECTED_6080,
  SV2V_UNCONNECTED_6081,SV2V_UNCONNECTED_6082,SV2V_UNCONNECTED_6083,
  SV2V_UNCONNECTED_6084,SV2V_UNCONNECTED_6085,SV2V_UNCONNECTED_6086,
  SV2V_UNCONNECTED_6087,SV2V_UNCONNECTED_6088,SV2V_UNCONNECTED_6089,
  SV2V_UNCONNECTED_6090,SV2V_UNCONNECTED_6091,SV2V_UNCONNECTED_6092,
  SV2V_UNCONNECTED_6093,SV2V_UNCONNECTED_6094,SV2V_UNCONNECTED_6095,
  SV2V_UNCONNECTED_6096,SV2V_UNCONNECTED_6097,SV2V_UNCONNECTED_6098,
  SV2V_UNCONNECTED_6099,SV2V_UNCONNECTED_6100,SV2V_UNCONNECTED_6101,
  SV2V_UNCONNECTED_6102,SV2V_UNCONNECTED_6103,SV2V_UNCONNECTED_6104,
  SV2V_UNCONNECTED_6105,SV2V_UNCONNECTED_6106,SV2V_UNCONNECTED_6107,SV2V_UNCONNECTED_6108,
  SV2V_UNCONNECTED_6109,SV2V_UNCONNECTED_6110,SV2V_UNCONNECTED_6111,
  SV2V_UNCONNECTED_6112,SV2V_UNCONNECTED_6113,SV2V_UNCONNECTED_6114,
  SV2V_UNCONNECTED_6115,SV2V_UNCONNECTED_6116,SV2V_UNCONNECTED_6117,
  SV2V_UNCONNECTED_6118,SV2V_UNCONNECTED_6119,SV2V_UNCONNECTED_6120,
  SV2V_UNCONNECTED_6121,SV2V_UNCONNECTED_6122,SV2V_UNCONNECTED_6123,
  SV2V_UNCONNECTED_6124,SV2V_UNCONNECTED_6125,SV2V_UNCONNECTED_6126,
  SV2V_UNCONNECTED_6127,SV2V_UNCONNECTED_6128,SV2V_UNCONNECTED_6129,
  SV2V_UNCONNECTED_6130,SV2V_UNCONNECTED_6131,SV2V_UNCONNECTED_6132,
  SV2V_UNCONNECTED_6133,SV2V_UNCONNECTED_6134,SV2V_UNCONNECTED_6135,
  SV2V_UNCONNECTED_6136,SV2V_UNCONNECTED_6137,SV2V_UNCONNECTED_6138,
  SV2V_UNCONNECTED_6139,SV2V_UNCONNECTED_6140,SV2V_UNCONNECTED_6141,
  SV2V_UNCONNECTED_6142,SV2V_UNCONNECTED_6143,SV2V_UNCONNECTED_6144,
  SV2V_UNCONNECTED_6145,SV2V_UNCONNECTED_6146,SV2V_UNCONNECTED_6147,SV2V_UNCONNECTED_6148,
  SV2V_UNCONNECTED_6149,SV2V_UNCONNECTED_6150,SV2V_UNCONNECTED_6151,
  SV2V_UNCONNECTED_6152,SV2V_UNCONNECTED_6153,SV2V_UNCONNECTED_6154,
  SV2V_UNCONNECTED_6155,SV2V_UNCONNECTED_6156,SV2V_UNCONNECTED_6157,
  SV2V_UNCONNECTED_6158,SV2V_UNCONNECTED_6159,SV2V_UNCONNECTED_6160,
  SV2V_UNCONNECTED_6161,SV2V_UNCONNECTED_6162,SV2V_UNCONNECTED_6163,
  SV2V_UNCONNECTED_6164,SV2V_UNCONNECTED_6165,SV2V_UNCONNECTED_6166,
  SV2V_UNCONNECTED_6167,SV2V_UNCONNECTED_6168,SV2V_UNCONNECTED_6169,
  SV2V_UNCONNECTED_6170,SV2V_UNCONNECTED_6171,SV2V_UNCONNECTED_6172,
  SV2V_UNCONNECTED_6173,SV2V_UNCONNECTED_6174,SV2V_UNCONNECTED_6175,
  SV2V_UNCONNECTED_6176,SV2V_UNCONNECTED_6177,SV2V_UNCONNECTED_6178,
  SV2V_UNCONNECTED_6179,SV2V_UNCONNECTED_6180,SV2V_UNCONNECTED_6181,
  SV2V_UNCONNECTED_6182,SV2V_UNCONNECTED_6183,SV2V_UNCONNECTED_6184,
  SV2V_UNCONNECTED_6185,SV2V_UNCONNECTED_6186,SV2V_UNCONNECTED_6187,SV2V_UNCONNECTED_6188,
  SV2V_UNCONNECTED_6189,SV2V_UNCONNECTED_6190,SV2V_UNCONNECTED_6191,
  SV2V_UNCONNECTED_6192,SV2V_UNCONNECTED_6193,SV2V_UNCONNECTED_6194,
  SV2V_UNCONNECTED_6195,SV2V_UNCONNECTED_6196,SV2V_UNCONNECTED_6197,
  SV2V_UNCONNECTED_6198,SV2V_UNCONNECTED_6199,SV2V_UNCONNECTED_6200,
  SV2V_UNCONNECTED_6201,SV2V_UNCONNECTED_6202,SV2V_UNCONNECTED_6203,
  SV2V_UNCONNECTED_6204,SV2V_UNCONNECTED_6205,SV2V_UNCONNECTED_6206,
  SV2V_UNCONNECTED_6207,SV2V_UNCONNECTED_6208,SV2V_UNCONNECTED_6209,
  SV2V_UNCONNECTED_6210,SV2V_UNCONNECTED_6211,SV2V_UNCONNECTED_6212,
  SV2V_UNCONNECTED_6213,SV2V_UNCONNECTED_6214,SV2V_UNCONNECTED_6215,
  SV2V_UNCONNECTED_6216,SV2V_UNCONNECTED_6217,SV2V_UNCONNECTED_6218,
  SV2V_UNCONNECTED_6219,SV2V_UNCONNECTED_6220,SV2V_UNCONNECTED_6221,
  SV2V_UNCONNECTED_6222,SV2V_UNCONNECTED_6223,SV2V_UNCONNECTED_6224,
  SV2V_UNCONNECTED_6225,SV2V_UNCONNECTED_6226,SV2V_UNCONNECTED_6227,SV2V_UNCONNECTED_6228,
  SV2V_UNCONNECTED_6229,SV2V_UNCONNECTED_6230,SV2V_UNCONNECTED_6231,
  SV2V_UNCONNECTED_6232,SV2V_UNCONNECTED_6233,SV2V_UNCONNECTED_6234,
  SV2V_UNCONNECTED_6235,SV2V_UNCONNECTED_6236,SV2V_UNCONNECTED_6237,
  SV2V_UNCONNECTED_6238,SV2V_UNCONNECTED_6239,SV2V_UNCONNECTED_6240,
  SV2V_UNCONNECTED_6241,SV2V_UNCONNECTED_6242,SV2V_UNCONNECTED_6243,
  SV2V_UNCONNECTED_6244,SV2V_UNCONNECTED_6245,SV2V_UNCONNECTED_6246,
  SV2V_UNCONNECTED_6247,SV2V_UNCONNECTED_6248,SV2V_UNCONNECTED_6249,
  SV2V_UNCONNECTED_6250,SV2V_UNCONNECTED_6251,SV2V_UNCONNECTED_6252,
  SV2V_UNCONNECTED_6253,SV2V_UNCONNECTED_6254,SV2V_UNCONNECTED_6255,
  SV2V_UNCONNECTED_6256,SV2V_UNCONNECTED_6257,SV2V_UNCONNECTED_6258,
  SV2V_UNCONNECTED_6259,SV2V_UNCONNECTED_6260,SV2V_UNCONNECTED_6261,
  SV2V_UNCONNECTED_6262,SV2V_UNCONNECTED_6263,SV2V_UNCONNECTED_6264,
  SV2V_UNCONNECTED_6265,SV2V_UNCONNECTED_6266,SV2V_UNCONNECTED_6267,SV2V_UNCONNECTED_6268,
  SV2V_UNCONNECTED_6269,SV2V_UNCONNECTED_6270,SV2V_UNCONNECTED_6271,
  SV2V_UNCONNECTED_6272,SV2V_UNCONNECTED_6273,SV2V_UNCONNECTED_6274,
  SV2V_UNCONNECTED_6275,SV2V_UNCONNECTED_6276,SV2V_UNCONNECTED_6277,
  SV2V_UNCONNECTED_6278,SV2V_UNCONNECTED_6279,SV2V_UNCONNECTED_6280,
  SV2V_UNCONNECTED_6281,SV2V_UNCONNECTED_6282,SV2V_UNCONNECTED_6283,
  SV2V_UNCONNECTED_6284,SV2V_UNCONNECTED_6285,SV2V_UNCONNECTED_6286,
  SV2V_UNCONNECTED_6287,SV2V_UNCONNECTED_6288,SV2V_UNCONNECTED_6289,
  SV2V_UNCONNECTED_6290,SV2V_UNCONNECTED_6291,SV2V_UNCONNECTED_6292,
  SV2V_UNCONNECTED_6293,SV2V_UNCONNECTED_6294,SV2V_UNCONNECTED_6295,
  SV2V_UNCONNECTED_6296,SV2V_UNCONNECTED_6297,SV2V_UNCONNECTED_6298,
  SV2V_UNCONNECTED_6299,SV2V_UNCONNECTED_6300,SV2V_UNCONNECTED_6301,
  SV2V_UNCONNECTED_6302,SV2V_UNCONNECTED_6303,SV2V_UNCONNECTED_6304,
  SV2V_UNCONNECTED_6305,SV2V_UNCONNECTED_6306,SV2V_UNCONNECTED_6307,SV2V_UNCONNECTED_6308,
  SV2V_UNCONNECTED_6309,SV2V_UNCONNECTED_6310,SV2V_UNCONNECTED_6311,
  SV2V_UNCONNECTED_6312,SV2V_UNCONNECTED_6313,SV2V_UNCONNECTED_6314,
  SV2V_UNCONNECTED_6315,SV2V_UNCONNECTED_6316,SV2V_UNCONNECTED_6317,
  SV2V_UNCONNECTED_6318,SV2V_UNCONNECTED_6319,SV2V_UNCONNECTED_6320,
  SV2V_UNCONNECTED_6321,SV2V_UNCONNECTED_6322,SV2V_UNCONNECTED_6323,
  SV2V_UNCONNECTED_6324,SV2V_UNCONNECTED_6325,SV2V_UNCONNECTED_6326,
  SV2V_UNCONNECTED_6327,SV2V_UNCONNECTED_6328,SV2V_UNCONNECTED_6329,
  SV2V_UNCONNECTED_6330,SV2V_UNCONNECTED_6331,SV2V_UNCONNECTED_6332,
  SV2V_UNCONNECTED_6333,SV2V_UNCONNECTED_6334,SV2V_UNCONNECTED_6335,
  SV2V_UNCONNECTED_6336,SV2V_UNCONNECTED_6337,SV2V_UNCONNECTED_6338,
  SV2V_UNCONNECTED_6339,SV2V_UNCONNECTED_6340,SV2V_UNCONNECTED_6341,
  SV2V_UNCONNECTED_6342,SV2V_UNCONNECTED_6343,SV2V_UNCONNECTED_6344,
  SV2V_UNCONNECTED_6345,SV2V_UNCONNECTED_6346,SV2V_UNCONNECTED_6347,SV2V_UNCONNECTED_6348,
  SV2V_UNCONNECTED_6349,SV2V_UNCONNECTED_6350,SV2V_UNCONNECTED_6351,
  SV2V_UNCONNECTED_6352,SV2V_UNCONNECTED_6353,SV2V_UNCONNECTED_6354,
  SV2V_UNCONNECTED_6355,SV2V_UNCONNECTED_6356,SV2V_UNCONNECTED_6357,
  SV2V_UNCONNECTED_6358,SV2V_UNCONNECTED_6359,SV2V_UNCONNECTED_6360,
  SV2V_UNCONNECTED_6361,SV2V_UNCONNECTED_6362,SV2V_UNCONNECTED_6363,
  SV2V_UNCONNECTED_6364,SV2V_UNCONNECTED_6365,SV2V_UNCONNECTED_6366,
  SV2V_UNCONNECTED_6367,SV2V_UNCONNECTED_6368,SV2V_UNCONNECTED_6369,
  SV2V_UNCONNECTED_6370,SV2V_UNCONNECTED_6371,SV2V_UNCONNECTED_6372,
  SV2V_UNCONNECTED_6373,SV2V_UNCONNECTED_6374,SV2V_UNCONNECTED_6375,
  SV2V_UNCONNECTED_6376,SV2V_UNCONNECTED_6377,SV2V_UNCONNECTED_6378,
  SV2V_UNCONNECTED_6379,SV2V_UNCONNECTED_6380,SV2V_UNCONNECTED_6381,
  SV2V_UNCONNECTED_6382,SV2V_UNCONNECTED_6383,SV2V_UNCONNECTED_6384,
  SV2V_UNCONNECTED_6385,SV2V_UNCONNECTED_6386,SV2V_UNCONNECTED_6387,SV2V_UNCONNECTED_6388,
  SV2V_UNCONNECTED_6389,SV2V_UNCONNECTED_6390,SV2V_UNCONNECTED_6391,
  SV2V_UNCONNECTED_6392,SV2V_UNCONNECTED_6393,SV2V_UNCONNECTED_6394,
  SV2V_UNCONNECTED_6395,SV2V_UNCONNECTED_6396,SV2V_UNCONNECTED_6397,
  SV2V_UNCONNECTED_6398,SV2V_UNCONNECTED_6399,SV2V_UNCONNECTED_6400,
  SV2V_UNCONNECTED_6401,SV2V_UNCONNECTED_6402,SV2V_UNCONNECTED_6403,
  SV2V_UNCONNECTED_6404,SV2V_UNCONNECTED_6405,SV2V_UNCONNECTED_6406,
  SV2V_UNCONNECTED_6407,SV2V_UNCONNECTED_6408,SV2V_UNCONNECTED_6409,
  SV2V_UNCONNECTED_6410,SV2V_UNCONNECTED_6411,SV2V_UNCONNECTED_6412,
  SV2V_UNCONNECTED_6413,SV2V_UNCONNECTED_6414,SV2V_UNCONNECTED_6415,
  SV2V_UNCONNECTED_6416,SV2V_UNCONNECTED_6417,SV2V_UNCONNECTED_6418,
  SV2V_UNCONNECTED_6419,SV2V_UNCONNECTED_6420,SV2V_UNCONNECTED_6421,
  SV2V_UNCONNECTED_6422,SV2V_UNCONNECTED_6423,SV2V_UNCONNECTED_6424,
  SV2V_UNCONNECTED_6425,SV2V_UNCONNECTED_6426,SV2V_UNCONNECTED_6427,SV2V_UNCONNECTED_6428,
  SV2V_UNCONNECTED_6429,SV2V_UNCONNECTED_6430,SV2V_UNCONNECTED_6431,
  SV2V_UNCONNECTED_6432,SV2V_UNCONNECTED_6433,SV2V_UNCONNECTED_6434,
  SV2V_UNCONNECTED_6435,SV2V_UNCONNECTED_6436,SV2V_UNCONNECTED_6437,
  SV2V_UNCONNECTED_6438,SV2V_UNCONNECTED_6439,SV2V_UNCONNECTED_6440,
  SV2V_UNCONNECTED_6441,SV2V_UNCONNECTED_6442,SV2V_UNCONNECTED_6443,
  SV2V_UNCONNECTED_6444,SV2V_UNCONNECTED_6445,SV2V_UNCONNECTED_6446,
  SV2V_UNCONNECTED_6447,SV2V_UNCONNECTED_6448,SV2V_UNCONNECTED_6449,
  SV2V_UNCONNECTED_6450,SV2V_UNCONNECTED_6451,SV2V_UNCONNECTED_6452,
  SV2V_UNCONNECTED_6453,SV2V_UNCONNECTED_6454,SV2V_UNCONNECTED_6455,
  SV2V_UNCONNECTED_6456,SV2V_UNCONNECTED_6457,SV2V_UNCONNECTED_6458,
  SV2V_UNCONNECTED_6459,SV2V_UNCONNECTED_6460,SV2V_UNCONNECTED_6461,
  SV2V_UNCONNECTED_6462,SV2V_UNCONNECTED_6463,SV2V_UNCONNECTED_6464,
  SV2V_UNCONNECTED_6465,SV2V_UNCONNECTED_6466,SV2V_UNCONNECTED_6467,SV2V_UNCONNECTED_6468,
  SV2V_UNCONNECTED_6469,SV2V_UNCONNECTED_6470,SV2V_UNCONNECTED_6471,
  SV2V_UNCONNECTED_6472,SV2V_UNCONNECTED_6473,SV2V_UNCONNECTED_6474,
  SV2V_UNCONNECTED_6475,SV2V_UNCONNECTED_6476,SV2V_UNCONNECTED_6477,
  SV2V_UNCONNECTED_6478,SV2V_UNCONNECTED_6479,SV2V_UNCONNECTED_6480,
  SV2V_UNCONNECTED_6481,SV2V_UNCONNECTED_6482,SV2V_UNCONNECTED_6483,
  SV2V_UNCONNECTED_6484,SV2V_UNCONNECTED_6485,SV2V_UNCONNECTED_6486,
  SV2V_UNCONNECTED_6487,SV2V_UNCONNECTED_6488,SV2V_UNCONNECTED_6489,
  SV2V_UNCONNECTED_6490,SV2V_UNCONNECTED_6491,SV2V_UNCONNECTED_6492,
  SV2V_UNCONNECTED_6493,SV2V_UNCONNECTED_6494,SV2V_UNCONNECTED_6495,
  SV2V_UNCONNECTED_6496,SV2V_UNCONNECTED_6497,SV2V_UNCONNECTED_6498,
  SV2V_UNCONNECTED_6499,SV2V_UNCONNECTED_6500,SV2V_UNCONNECTED_6501,
  SV2V_UNCONNECTED_6502,SV2V_UNCONNECTED_6503,SV2V_UNCONNECTED_6504,
  SV2V_UNCONNECTED_6505,SV2V_UNCONNECTED_6506,SV2V_UNCONNECTED_6507,SV2V_UNCONNECTED_6508,
  SV2V_UNCONNECTED_6509,SV2V_UNCONNECTED_6510,SV2V_UNCONNECTED_6511,
  SV2V_UNCONNECTED_6512,SV2V_UNCONNECTED_6513,SV2V_UNCONNECTED_6514,
  SV2V_UNCONNECTED_6515,SV2V_UNCONNECTED_6516,SV2V_UNCONNECTED_6517,
  SV2V_UNCONNECTED_6518,SV2V_UNCONNECTED_6519,SV2V_UNCONNECTED_6520,
  SV2V_UNCONNECTED_6521,SV2V_UNCONNECTED_6522,SV2V_UNCONNECTED_6523,
  SV2V_UNCONNECTED_6524,SV2V_UNCONNECTED_6525,SV2V_UNCONNECTED_6526,
  SV2V_UNCONNECTED_6527,SV2V_UNCONNECTED_6528,SV2V_UNCONNECTED_6529,
  SV2V_UNCONNECTED_6530,SV2V_UNCONNECTED_6531,SV2V_UNCONNECTED_6532,
  SV2V_UNCONNECTED_6533,SV2V_UNCONNECTED_6534,SV2V_UNCONNECTED_6535,
  SV2V_UNCONNECTED_6536,SV2V_UNCONNECTED_6537,SV2V_UNCONNECTED_6538,
  SV2V_UNCONNECTED_6539,SV2V_UNCONNECTED_6540,SV2V_UNCONNECTED_6541,
  SV2V_UNCONNECTED_6542,SV2V_UNCONNECTED_6543,SV2V_UNCONNECTED_6544,
  SV2V_UNCONNECTED_6545,SV2V_UNCONNECTED_6546,SV2V_UNCONNECTED_6547,SV2V_UNCONNECTED_6548,
  SV2V_UNCONNECTED_6549,SV2V_UNCONNECTED_6550,SV2V_UNCONNECTED_6551,
  SV2V_UNCONNECTED_6552,SV2V_UNCONNECTED_6553,SV2V_UNCONNECTED_6554,
  SV2V_UNCONNECTED_6555,SV2V_UNCONNECTED_6556,SV2V_UNCONNECTED_6557,
  SV2V_UNCONNECTED_6558,SV2V_UNCONNECTED_6559,SV2V_UNCONNECTED_6560,
  SV2V_UNCONNECTED_6561,SV2V_UNCONNECTED_6562,SV2V_UNCONNECTED_6563,
  SV2V_UNCONNECTED_6564,SV2V_UNCONNECTED_6565,SV2V_UNCONNECTED_6566,
  SV2V_UNCONNECTED_6567,SV2V_UNCONNECTED_6568,SV2V_UNCONNECTED_6569,
  SV2V_UNCONNECTED_6570,SV2V_UNCONNECTED_6571,SV2V_UNCONNECTED_6572,
  SV2V_UNCONNECTED_6573,SV2V_UNCONNECTED_6574,SV2V_UNCONNECTED_6575,
  SV2V_UNCONNECTED_6576,SV2V_UNCONNECTED_6577,SV2V_UNCONNECTED_6578,
  SV2V_UNCONNECTED_6579,SV2V_UNCONNECTED_6580,SV2V_UNCONNECTED_6581,
  SV2V_UNCONNECTED_6582,SV2V_UNCONNECTED_6583,SV2V_UNCONNECTED_6584,
  SV2V_UNCONNECTED_6585,SV2V_UNCONNECTED_6586,SV2V_UNCONNECTED_6587,SV2V_UNCONNECTED_6588,
  SV2V_UNCONNECTED_6589,SV2V_UNCONNECTED_6590,SV2V_UNCONNECTED_6591,
  SV2V_UNCONNECTED_6592,SV2V_UNCONNECTED_6593,SV2V_UNCONNECTED_6594,
  SV2V_UNCONNECTED_6595,SV2V_UNCONNECTED_6596,SV2V_UNCONNECTED_6597,
  SV2V_UNCONNECTED_6598,SV2V_UNCONNECTED_6599,SV2V_UNCONNECTED_6600,
  SV2V_UNCONNECTED_6601,SV2V_UNCONNECTED_6602,SV2V_UNCONNECTED_6603,
  SV2V_UNCONNECTED_6604,SV2V_UNCONNECTED_6605,SV2V_UNCONNECTED_6606,
  SV2V_UNCONNECTED_6607,SV2V_UNCONNECTED_6608,SV2V_UNCONNECTED_6609,
  SV2V_UNCONNECTED_6610,SV2V_UNCONNECTED_6611,SV2V_UNCONNECTED_6612,
  SV2V_UNCONNECTED_6613,SV2V_UNCONNECTED_6614,SV2V_UNCONNECTED_6615,
  SV2V_UNCONNECTED_6616,SV2V_UNCONNECTED_6617,SV2V_UNCONNECTED_6618,
  SV2V_UNCONNECTED_6619,SV2V_UNCONNECTED_6620,SV2V_UNCONNECTED_6621,
  SV2V_UNCONNECTED_6622,SV2V_UNCONNECTED_6623,SV2V_UNCONNECTED_6624,
  SV2V_UNCONNECTED_6625,SV2V_UNCONNECTED_6626,SV2V_UNCONNECTED_6627,SV2V_UNCONNECTED_6628,
  SV2V_UNCONNECTED_6629,SV2V_UNCONNECTED_6630,SV2V_UNCONNECTED_6631,
  SV2V_UNCONNECTED_6632,SV2V_UNCONNECTED_6633,SV2V_UNCONNECTED_6634,
  SV2V_UNCONNECTED_6635,SV2V_UNCONNECTED_6636,SV2V_UNCONNECTED_6637,
  SV2V_UNCONNECTED_6638,SV2V_UNCONNECTED_6639,SV2V_UNCONNECTED_6640,
  SV2V_UNCONNECTED_6641,SV2V_UNCONNECTED_6642,SV2V_UNCONNECTED_6643,
  SV2V_UNCONNECTED_6644,SV2V_UNCONNECTED_6645,SV2V_UNCONNECTED_6646,
  SV2V_UNCONNECTED_6647,SV2V_UNCONNECTED_6648,SV2V_UNCONNECTED_6649,
  SV2V_UNCONNECTED_6650,SV2V_UNCONNECTED_6651,SV2V_UNCONNECTED_6652,
  SV2V_UNCONNECTED_6653,SV2V_UNCONNECTED_6654,SV2V_UNCONNECTED_6655,
  SV2V_UNCONNECTED_6656,SV2V_UNCONNECTED_6657,SV2V_UNCONNECTED_6658,
  SV2V_UNCONNECTED_6659,SV2V_UNCONNECTED_6660,SV2V_UNCONNECTED_6661,
  SV2V_UNCONNECTED_6662,SV2V_UNCONNECTED_6663,SV2V_UNCONNECTED_6664,
  SV2V_UNCONNECTED_6665,SV2V_UNCONNECTED_6666,SV2V_UNCONNECTED_6667,SV2V_UNCONNECTED_6668,
  SV2V_UNCONNECTED_6669,SV2V_UNCONNECTED_6670,SV2V_UNCONNECTED_6671,
  SV2V_UNCONNECTED_6672,SV2V_UNCONNECTED_6673,SV2V_UNCONNECTED_6674,
  SV2V_UNCONNECTED_6675,SV2V_UNCONNECTED_6676,SV2V_UNCONNECTED_6677,
  SV2V_UNCONNECTED_6678,SV2V_UNCONNECTED_6679,SV2V_UNCONNECTED_6680,
  SV2V_UNCONNECTED_6681,SV2V_UNCONNECTED_6682,SV2V_UNCONNECTED_6683,
  SV2V_UNCONNECTED_6684,SV2V_UNCONNECTED_6685,SV2V_UNCONNECTED_6686,
  SV2V_UNCONNECTED_6687,SV2V_UNCONNECTED_6688,SV2V_UNCONNECTED_6689,
  SV2V_UNCONNECTED_6690,SV2V_UNCONNECTED_6691,SV2V_UNCONNECTED_6692,
  SV2V_UNCONNECTED_6693,SV2V_UNCONNECTED_6694,SV2V_UNCONNECTED_6695,
  SV2V_UNCONNECTED_6696,SV2V_UNCONNECTED_6697,SV2V_UNCONNECTED_6698,
  SV2V_UNCONNECTED_6699,SV2V_UNCONNECTED_6700,SV2V_UNCONNECTED_6701,
  SV2V_UNCONNECTED_6702,SV2V_UNCONNECTED_6703,SV2V_UNCONNECTED_6704,
  SV2V_UNCONNECTED_6705,SV2V_UNCONNECTED_6706,SV2V_UNCONNECTED_6707,SV2V_UNCONNECTED_6708,
  SV2V_UNCONNECTED_6709,SV2V_UNCONNECTED_6710,SV2V_UNCONNECTED_6711,
  SV2V_UNCONNECTED_6712,SV2V_UNCONNECTED_6713,SV2V_UNCONNECTED_6714,
  SV2V_UNCONNECTED_6715,SV2V_UNCONNECTED_6716,SV2V_UNCONNECTED_6717,
  SV2V_UNCONNECTED_6718,SV2V_UNCONNECTED_6719,SV2V_UNCONNECTED_6720,
  SV2V_UNCONNECTED_6721,SV2V_UNCONNECTED_6722,SV2V_UNCONNECTED_6723,
  SV2V_UNCONNECTED_6724,SV2V_UNCONNECTED_6725,SV2V_UNCONNECTED_6726,
  SV2V_UNCONNECTED_6727,SV2V_UNCONNECTED_6728,SV2V_UNCONNECTED_6729,
  SV2V_UNCONNECTED_6730,SV2V_UNCONNECTED_6731,SV2V_UNCONNECTED_6732,
  SV2V_UNCONNECTED_6733,SV2V_UNCONNECTED_6734,SV2V_UNCONNECTED_6735,
  SV2V_UNCONNECTED_6736,SV2V_UNCONNECTED_6737,SV2V_UNCONNECTED_6738,
  SV2V_UNCONNECTED_6739,SV2V_UNCONNECTED_6740,SV2V_UNCONNECTED_6741,
  SV2V_UNCONNECTED_6742,SV2V_UNCONNECTED_6743,SV2V_UNCONNECTED_6744,
  SV2V_UNCONNECTED_6745,SV2V_UNCONNECTED_6746,SV2V_UNCONNECTED_6747,SV2V_UNCONNECTED_6748,
  SV2V_UNCONNECTED_6749,SV2V_UNCONNECTED_6750,SV2V_UNCONNECTED_6751,
  SV2V_UNCONNECTED_6752,SV2V_UNCONNECTED_6753,SV2V_UNCONNECTED_6754,
  SV2V_UNCONNECTED_6755,SV2V_UNCONNECTED_6756,SV2V_UNCONNECTED_6757,
  SV2V_UNCONNECTED_6758,SV2V_UNCONNECTED_6759,SV2V_UNCONNECTED_6760,
  SV2V_UNCONNECTED_6761,SV2V_UNCONNECTED_6762,SV2V_UNCONNECTED_6763,
  SV2V_UNCONNECTED_6764,SV2V_UNCONNECTED_6765,SV2V_UNCONNECTED_6766,
  SV2V_UNCONNECTED_6767,SV2V_UNCONNECTED_6768,SV2V_UNCONNECTED_6769,
  SV2V_UNCONNECTED_6770,SV2V_UNCONNECTED_6771,SV2V_UNCONNECTED_6772,
  SV2V_UNCONNECTED_6773,SV2V_UNCONNECTED_6774,SV2V_UNCONNECTED_6775,
  SV2V_UNCONNECTED_6776,SV2V_UNCONNECTED_6777,SV2V_UNCONNECTED_6778,
  SV2V_UNCONNECTED_6779,SV2V_UNCONNECTED_6780,SV2V_UNCONNECTED_6781,
  SV2V_UNCONNECTED_6782,SV2V_UNCONNECTED_6783,SV2V_UNCONNECTED_6784,
  SV2V_UNCONNECTED_6785,SV2V_UNCONNECTED_6786,SV2V_UNCONNECTED_6787,SV2V_UNCONNECTED_6788,
  SV2V_UNCONNECTED_6789,SV2V_UNCONNECTED_6790,SV2V_UNCONNECTED_6791,
  SV2V_UNCONNECTED_6792,SV2V_UNCONNECTED_6793,SV2V_UNCONNECTED_6794,
  SV2V_UNCONNECTED_6795,SV2V_UNCONNECTED_6796,SV2V_UNCONNECTED_6797,
  SV2V_UNCONNECTED_6798,SV2V_UNCONNECTED_6799,SV2V_UNCONNECTED_6800,
  SV2V_UNCONNECTED_6801,SV2V_UNCONNECTED_6802,SV2V_UNCONNECTED_6803,
  SV2V_UNCONNECTED_6804,SV2V_UNCONNECTED_6805,SV2V_UNCONNECTED_6806,
  SV2V_UNCONNECTED_6807,SV2V_UNCONNECTED_6808,SV2V_UNCONNECTED_6809,
  SV2V_UNCONNECTED_6810,SV2V_UNCONNECTED_6811,SV2V_UNCONNECTED_6812,
  SV2V_UNCONNECTED_6813,SV2V_UNCONNECTED_6814,SV2V_UNCONNECTED_6815,
  SV2V_UNCONNECTED_6816,SV2V_UNCONNECTED_6817,SV2V_UNCONNECTED_6818,
  SV2V_UNCONNECTED_6819,SV2V_UNCONNECTED_6820,SV2V_UNCONNECTED_6821,
  SV2V_UNCONNECTED_6822,SV2V_UNCONNECTED_6823,SV2V_UNCONNECTED_6824,
  SV2V_UNCONNECTED_6825,SV2V_UNCONNECTED_6826,SV2V_UNCONNECTED_6827,SV2V_UNCONNECTED_6828,
  SV2V_UNCONNECTED_6829,SV2V_UNCONNECTED_6830,SV2V_UNCONNECTED_6831,
  SV2V_UNCONNECTED_6832,SV2V_UNCONNECTED_6833,SV2V_UNCONNECTED_6834,
  SV2V_UNCONNECTED_6835,SV2V_UNCONNECTED_6836,SV2V_UNCONNECTED_6837,
  SV2V_UNCONNECTED_6838,SV2V_UNCONNECTED_6839,SV2V_UNCONNECTED_6840,
  SV2V_UNCONNECTED_6841,SV2V_UNCONNECTED_6842,SV2V_UNCONNECTED_6843,
  SV2V_UNCONNECTED_6844,SV2V_UNCONNECTED_6845,SV2V_UNCONNECTED_6846,
  SV2V_UNCONNECTED_6847,SV2V_UNCONNECTED_6848,SV2V_UNCONNECTED_6849,
  SV2V_UNCONNECTED_6850,SV2V_UNCONNECTED_6851,SV2V_UNCONNECTED_6852,
  SV2V_UNCONNECTED_6853,SV2V_UNCONNECTED_6854,SV2V_UNCONNECTED_6855,
  SV2V_UNCONNECTED_6856,SV2V_UNCONNECTED_6857,SV2V_UNCONNECTED_6858,
  SV2V_UNCONNECTED_6859,SV2V_UNCONNECTED_6860,SV2V_UNCONNECTED_6861,
  SV2V_UNCONNECTED_6862,SV2V_UNCONNECTED_6863,SV2V_UNCONNECTED_6864,
  SV2V_UNCONNECTED_6865,SV2V_UNCONNECTED_6866,SV2V_UNCONNECTED_6867,SV2V_UNCONNECTED_6868,
  SV2V_UNCONNECTED_6869,SV2V_UNCONNECTED_6870,SV2V_UNCONNECTED_6871,
  SV2V_UNCONNECTED_6872,SV2V_UNCONNECTED_6873,SV2V_UNCONNECTED_6874,
  SV2V_UNCONNECTED_6875,SV2V_UNCONNECTED_6876,SV2V_UNCONNECTED_6877,
  SV2V_UNCONNECTED_6878,SV2V_UNCONNECTED_6879,SV2V_UNCONNECTED_6880,
  SV2V_UNCONNECTED_6881,SV2V_UNCONNECTED_6882,SV2V_UNCONNECTED_6883,
  SV2V_UNCONNECTED_6884,SV2V_UNCONNECTED_6885,SV2V_UNCONNECTED_6886,
  SV2V_UNCONNECTED_6887,SV2V_UNCONNECTED_6888,SV2V_UNCONNECTED_6889,
  SV2V_UNCONNECTED_6890,SV2V_UNCONNECTED_6891,SV2V_UNCONNECTED_6892,
  SV2V_UNCONNECTED_6893,SV2V_UNCONNECTED_6894,SV2V_UNCONNECTED_6895,
  SV2V_UNCONNECTED_6896,SV2V_UNCONNECTED_6897,SV2V_UNCONNECTED_6898,
  SV2V_UNCONNECTED_6899,SV2V_UNCONNECTED_6900,SV2V_UNCONNECTED_6901,
  SV2V_UNCONNECTED_6902,SV2V_UNCONNECTED_6903,SV2V_UNCONNECTED_6904,
  SV2V_UNCONNECTED_6905,SV2V_UNCONNECTED_6906,SV2V_UNCONNECTED_6907,SV2V_UNCONNECTED_6908,
  SV2V_UNCONNECTED_6909,SV2V_UNCONNECTED_6910,SV2V_UNCONNECTED_6911,
  SV2V_UNCONNECTED_6912,SV2V_UNCONNECTED_6913,SV2V_UNCONNECTED_6914,
  SV2V_UNCONNECTED_6915,SV2V_UNCONNECTED_6916,SV2V_UNCONNECTED_6917,
  SV2V_UNCONNECTED_6918,SV2V_UNCONNECTED_6919,SV2V_UNCONNECTED_6920,
  SV2V_UNCONNECTED_6921,SV2V_UNCONNECTED_6922,SV2V_UNCONNECTED_6923,
  SV2V_UNCONNECTED_6924,SV2V_UNCONNECTED_6925,SV2V_UNCONNECTED_6926,
  SV2V_UNCONNECTED_6927,SV2V_UNCONNECTED_6928,SV2V_UNCONNECTED_6929,
  SV2V_UNCONNECTED_6930,SV2V_UNCONNECTED_6931,SV2V_UNCONNECTED_6932,
  SV2V_UNCONNECTED_6933,SV2V_UNCONNECTED_6934,SV2V_UNCONNECTED_6935,
  SV2V_UNCONNECTED_6936,SV2V_UNCONNECTED_6937,SV2V_UNCONNECTED_6938,
  SV2V_UNCONNECTED_6939,SV2V_UNCONNECTED_6940,SV2V_UNCONNECTED_6941,
  SV2V_UNCONNECTED_6942,SV2V_UNCONNECTED_6943,SV2V_UNCONNECTED_6944,
  SV2V_UNCONNECTED_6945,SV2V_UNCONNECTED_6946,SV2V_UNCONNECTED_6947,SV2V_UNCONNECTED_6948,
  SV2V_UNCONNECTED_6949,SV2V_UNCONNECTED_6950,SV2V_UNCONNECTED_6951,
  SV2V_UNCONNECTED_6952,SV2V_UNCONNECTED_6953,SV2V_UNCONNECTED_6954,
  SV2V_UNCONNECTED_6955,SV2V_UNCONNECTED_6956,SV2V_UNCONNECTED_6957,
  SV2V_UNCONNECTED_6958,SV2V_UNCONNECTED_6959,SV2V_UNCONNECTED_6960,
  SV2V_UNCONNECTED_6961,SV2V_UNCONNECTED_6962,SV2V_UNCONNECTED_6963,
  SV2V_UNCONNECTED_6964,SV2V_UNCONNECTED_6965,SV2V_UNCONNECTED_6966,
  SV2V_UNCONNECTED_6967,SV2V_UNCONNECTED_6968,SV2V_UNCONNECTED_6969,
  SV2V_UNCONNECTED_6970,SV2V_UNCONNECTED_6971,SV2V_UNCONNECTED_6972,
  SV2V_UNCONNECTED_6973,SV2V_UNCONNECTED_6974,SV2V_UNCONNECTED_6975,
  SV2V_UNCONNECTED_6976,SV2V_UNCONNECTED_6977,SV2V_UNCONNECTED_6978,
  SV2V_UNCONNECTED_6979,SV2V_UNCONNECTED_6980,SV2V_UNCONNECTED_6981,
  SV2V_UNCONNECTED_6982,SV2V_UNCONNECTED_6983,SV2V_UNCONNECTED_6984,
  SV2V_UNCONNECTED_6985,SV2V_UNCONNECTED_6986,SV2V_UNCONNECTED_6987,SV2V_UNCONNECTED_6988,
  SV2V_UNCONNECTED_6989,SV2V_UNCONNECTED_6990,SV2V_UNCONNECTED_6991,
  SV2V_UNCONNECTED_6992,SV2V_UNCONNECTED_6993,SV2V_UNCONNECTED_6994,
  SV2V_UNCONNECTED_6995,SV2V_UNCONNECTED_6996,SV2V_UNCONNECTED_6997,
  SV2V_UNCONNECTED_6998,SV2V_UNCONNECTED_6999,SV2V_UNCONNECTED_7000,
  SV2V_UNCONNECTED_7001,SV2V_UNCONNECTED_7002,SV2V_UNCONNECTED_7003,
  SV2V_UNCONNECTED_7004,SV2V_UNCONNECTED_7005,SV2V_UNCONNECTED_7006,
  SV2V_UNCONNECTED_7007,SV2V_UNCONNECTED_7008,SV2V_UNCONNECTED_7009,
  SV2V_UNCONNECTED_7010,SV2V_UNCONNECTED_7011,SV2V_UNCONNECTED_7012,
  SV2V_UNCONNECTED_7013,SV2V_UNCONNECTED_7014,SV2V_UNCONNECTED_7015,
  SV2V_UNCONNECTED_7016,SV2V_UNCONNECTED_7017,SV2V_UNCONNECTED_7018,
  SV2V_UNCONNECTED_7019,SV2V_UNCONNECTED_7020,SV2V_UNCONNECTED_7021,
  SV2V_UNCONNECTED_7022,SV2V_UNCONNECTED_7023,SV2V_UNCONNECTED_7024,
  SV2V_UNCONNECTED_7025,SV2V_UNCONNECTED_7026,SV2V_UNCONNECTED_7027,SV2V_UNCONNECTED_7028,
  SV2V_UNCONNECTED_7029,SV2V_UNCONNECTED_7030,SV2V_UNCONNECTED_7031,
  SV2V_UNCONNECTED_7032,SV2V_UNCONNECTED_7033,SV2V_UNCONNECTED_7034,
  SV2V_UNCONNECTED_7035,SV2V_UNCONNECTED_7036,SV2V_UNCONNECTED_7037,
  SV2V_UNCONNECTED_7038,SV2V_UNCONNECTED_7039,SV2V_UNCONNECTED_7040,
  SV2V_UNCONNECTED_7041,SV2V_UNCONNECTED_7042,SV2V_UNCONNECTED_7043,
  SV2V_UNCONNECTED_7044,SV2V_UNCONNECTED_7045,SV2V_UNCONNECTED_7046,
  SV2V_UNCONNECTED_7047,SV2V_UNCONNECTED_7048,SV2V_UNCONNECTED_7049,
  SV2V_UNCONNECTED_7050,SV2V_UNCONNECTED_7051,SV2V_UNCONNECTED_7052,
  SV2V_UNCONNECTED_7053,SV2V_UNCONNECTED_7054,SV2V_UNCONNECTED_7055,
  SV2V_UNCONNECTED_7056,SV2V_UNCONNECTED_7057,SV2V_UNCONNECTED_7058,
  SV2V_UNCONNECTED_7059,SV2V_UNCONNECTED_7060,SV2V_UNCONNECTED_7061,
  SV2V_UNCONNECTED_7062,SV2V_UNCONNECTED_7063,SV2V_UNCONNECTED_7064,
  SV2V_UNCONNECTED_7065,SV2V_UNCONNECTED_7066,SV2V_UNCONNECTED_7067,SV2V_UNCONNECTED_7068,
  SV2V_UNCONNECTED_7069,SV2V_UNCONNECTED_7070,SV2V_UNCONNECTED_7071,
  SV2V_UNCONNECTED_7072,SV2V_UNCONNECTED_7073,SV2V_UNCONNECTED_7074,
  SV2V_UNCONNECTED_7075,SV2V_UNCONNECTED_7076,SV2V_UNCONNECTED_7077,
  SV2V_UNCONNECTED_7078,SV2V_UNCONNECTED_7079,SV2V_UNCONNECTED_7080,
  SV2V_UNCONNECTED_7081,SV2V_UNCONNECTED_7082,SV2V_UNCONNECTED_7083,
  SV2V_UNCONNECTED_7084,SV2V_UNCONNECTED_7085,SV2V_UNCONNECTED_7086,
  SV2V_UNCONNECTED_7087,SV2V_UNCONNECTED_7088,SV2V_UNCONNECTED_7089,
  SV2V_UNCONNECTED_7090,SV2V_UNCONNECTED_7091,SV2V_UNCONNECTED_7092,
  SV2V_UNCONNECTED_7093,SV2V_UNCONNECTED_7094,SV2V_UNCONNECTED_7095,
  SV2V_UNCONNECTED_7096,SV2V_UNCONNECTED_7097,SV2V_UNCONNECTED_7098,
  SV2V_UNCONNECTED_7099,SV2V_UNCONNECTED_7100,SV2V_UNCONNECTED_7101,
  SV2V_UNCONNECTED_7102,SV2V_UNCONNECTED_7103,SV2V_UNCONNECTED_7104,
  SV2V_UNCONNECTED_7105,SV2V_UNCONNECTED_7106,SV2V_UNCONNECTED_7107,SV2V_UNCONNECTED_7108,
  SV2V_UNCONNECTED_7109,SV2V_UNCONNECTED_7110,SV2V_UNCONNECTED_7111,
  SV2V_UNCONNECTED_7112,SV2V_UNCONNECTED_7113,SV2V_UNCONNECTED_7114,
  SV2V_UNCONNECTED_7115,SV2V_UNCONNECTED_7116,SV2V_UNCONNECTED_7117,
  SV2V_UNCONNECTED_7118,SV2V_UNCONNECTED_7119,SV2V_UNCONNECTED_7120,
  SV2V_UNCONNECTED_7121,SV2V_UNCONNECTED_7122,SV2V_UNCONNECTED_7123,
  SV2V_UNCONNECTED_7124,SV2V_UNCONNECTED_7125,SV2V_UNCONNECTED_7126,
  SV2V_UNCONNECTED_7127,SV2V_UNCONNECTED_7128,SV2V_UNCONNECTED_7129,
  SV2V_UNCONNECTED_7130,SV2V_UNCONNECTED_7131,SV2V_UNCONNECTED_7132,
  SV2V_UNCONNECTED_7133,SV2V_UNCONNECTED_7134,SV2V_UNCONNECTED_7135,
  SV2V_UNCONNECTED_7136,SV2V_UNCONNECTED_7137,SV2V_UNCONNECTED_7138,
  SV2V_UNCONNECTED_7139,SV2V_UNCONNECTED_7140,SV2V_UNCONNECTED_7141,
  SV2V_UNCONNECTED_7142,SV2V_UNCONNECTED_7143,SV2V_UNCONNECTED_7144,
  SV2V_UNCONNECTED_7145,SV2V_UNCONNECTED_7146,SV2V_UNCONNECTED_7147,SV2V_UNCONNECTED_7148,
  SV2V_UNCONNECTED_7149,SV2V_UNCONNECTED_7150,SV2V_UNCONNECTED_7151,
  SV2V_UNCONNECTED_7152,SV2V_UNCONNECTED_7153,SV2V_UNCONNECTED_7154,
  SV2V_UNCONNECTED_7155,SV2V_UNCONNECTED_7156,SV2V_UNCONNECTED_7157,
  SV2V_UNCONNECTED_7158,SV2V_UNCONNECTED_7159,SV2V_UNCONNECTED_7160,
  SV2V_UNCONNECTED_7161,SV2V_UNCONNECTED_7162,SV2V_UNCONNECTED_7163,
  SV2V_UNCONNECTED_7164,SV2V_UNCONNECTED_7165,SV2V_UNCONNECTED_7166,
  SV2V_UNCONNECTED_7167;
  wire [55:54] T885,T2;
  wire [1:0] T169,T73,T720,T722;
  wire [1:1] T4,T891;
  wire [52:0] T9,T10,T899,T239,T242,T246,T927,T489,T488,T494,T499,T503,T505,T513,T506,T514,
  T581,T673,T700,T701;
  wire [2:0] T28,T29,T36,T38,T43,T45,T71,T72,T80,T84,T81,T82;
  wire [3:2] T78;
  wire [2:2] T85;
  wire [13:0] T196,T197,T594,T604,T595,expP1_PC,T759,T766,T760,T772,T767;
  wire [11:0] T198,T311,T315,T319,T323,T327,T331,T827,T832,T834,T837,T840,T838,T843,T841,T846,
  T844,T847;
  wire [53:53] T897;
  wire [104:47] T217,T233;
  wire [103:46] T898;
  wire [32:0] T900;
  wire [29:0] T901;
  wire [45:0] T902,T244,T930;
  wire [51:0] T925,sigY_E1,T724,T715,roundEvenMask_E1,sigY1_E,sigY0_E,T725,T816,T819;
  wire [52:36] T247,T516;
  wire [16:0] ER1_A1_sqrt;
  wire [14:0] T903;
  wire [15:0] T251,T587;
  wire [8:0] mulAdd9Out_A,T258,zFractR0_A6_sqrt,zFractR0_A4_div,T260,T265,mulAdd9A_A,
  mulAdd9B_A,T408,T388,T390,T394,T391,T397,T395,T398,T401,T399,T402,zK1_A4_div,T411,T413,
  T415,T417,T419,T421,T451,T424,T917,T426,T432,T919,T428,T436,T920,T438,T921,T441,
  T922,T442,T443,zK2_A7_sqrt,T453,T455;
  wire [18:18] loMulAdd9Out_A;
  wire [17:0] T916,T253;
  wire [24:18] mulAdd9C_A;
  wire [24:0] T271;
  wire [23:15] T904;
  wire [20:0] T905,T282,T275,T277,T295,T283,T284,T300,T304;
  wire [24:16] T272;
  wire [9:0] T292,T369,T375;
  wire [9:1] sqrR0_A5_sqrt;
  wire [10:10] T910,T328,T842;
  wire [19:0] T911,T302,T914;
  wire [20:7] T305;
  wire [11:11] T308,T312,T316,T320,T324,T353,T826,T828,T833,T845,T848;
  wire [4:4] T335,T358;
  wire [9:9] T332,T365,T835,T839;
  wire [19:10] T364;
  wire [18:5] T339;
  wire [12:0] T346,T352,T590,posExpX_E,T933,T592,T709,T943,T711;
  wire [12:12] T342,T347;
  wire [8:8] T370,T376,T420,T423,T422,T454,T457;
  wire [5:5] T381;
  wire [7:7] T410,T412,T414,T416,T418,T452,T456;
  wire [48:44] zFractB_A4_div;
  wire [6:0] T461;
  wire [51:36] T475;
  wire [50:19] T926;
  wire [45:15] T928;
  wire [45:13] T929;
  wire [51:4] T932;
  wire [0:0] roundMask_E,expP2_PC,incrPosMask_E,T944,T946;
  wire [31:0] T588;
  wire [13:13] sExpX_E,sExpY_E1;
  wire [13:1] T598;
  wire [15:15] T618,T621;
  wire [14:14] T619;
  wire [15:14] T622,T625;
  wire [13:12] T623;
  wire [15:12] T626,T629;
  wire [11:8] T627;
  wire [31:31] T643,T646;
  wire [30:30] T644;
  wire [31:30] T647,T650;
  wire [29:28] T648;
  wire [31:28] T651,T654;
  wire [27:24] T652;
  wire [31:24] T655,T658;
  wire [23:16] T656;
  wire [51:51] T812,T817;
  reg extraT_E,sqrtOp_PC,sqrtOp_PB,sqrtOp_PA,sign_PC,sign_PB,sign_PA,valid_PC,
  valid_PA,valid_PB,sigB_PA_50,sigB_PA_49,sigB_PA_48,sigB_PA_47,fractB_51_PB,sigB_PA_51,
  fractA_0_PB,E_E_div,sqrSigma1_C_0,isZeroRemT_E,isNegRemT_E,fractA_51_PC,
  fractA_51_PB;
  reg [2:0] cycleNum_E,cycleNum_C,cycleNum_A;
  reg [1:0] T51,T114,T137,T53,T116,T139,T170,roundingMode_PC,roundingMode_PB,
  roundingMode_PA;
  reg [0:0] specialCodeB_PC,specialCodeB_PB,specialCodeB_PA,specialCodeA_PC,specialCodeA_PB,
  specialCodeA_PA,exp_PC;
  reg [3:0] cycleNum_B;
  reg [51:1] sigB_PC;
  reg [50:0] fractB_other_PB;
  reg [20:0] T285,partNegSigma0_A;
  reg [25:0] sigB_PA;
  reg [12:0] T593;
  reg [13:0] exp_PB,exp_PA;
  reg [53:53] T206;
  reg [51:0] sigA_PA;
  reg [104:47] T218;
  reg [103:46] T230;
  reg [32:31] sqrSigma1_C;
  reg [29:0] T241;
  reg [52:36] T248;
  reg [23:15] T256;
  reg [9:0] T908;
  reg [8:0] nextMulAdd9B_A,T918;
  reg [50:19] T472;
  reg [45:15] T491;
  reg [52:0] T727;
  assign T707 = posExpX_E <= { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 };
  assign T708 = T709 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign T776 = { 1'b1, 1'b1 } <= T709[12:10];

  always @(posedge clk) begin
    if(N312) begin
      extraT_E <= sigT_C1[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      sqrtOp_PC <= T17;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      sqrtOp_PB <= T19;
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      sqrtOp_PA <= io_sqrtOp;
    end 
  end


  always @(posedge clk) begin
    if(N169) begin
      cycleNum_E[2] <= N172;
    end 
  end


  always @(posedge clk) begin
    if(N169) begin
      cycleNum_E[1] <= N171;
    end 
  end


  always @(posedge clk) begin
    if(N169) begin
      cycleNum_E[0] <= N170;
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      T51[1] <= T36[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      T51[0] <= T36[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      specialCodeB_PC[0] <= T36[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      T114[1] <= T38[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      T114[0] <= T38[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      specialCodeB_PB[0] <= T38[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      T137[1] <= io_b[63];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      T137[0] <= io_b[62];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      specialCodeB_PA[0] <= io_b[61];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      T53[1] <= T43[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      T53[0] <= T43[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      specialCodeA_PC[0] <= T43[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      T116[1] <= T45[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      T116[0] <= T45[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      specialCodeA_PB[0] <= T45[0];
    end 
  end


  always @(posedge clk) begin
    if(T47) begin
      T139[1] <= io_a[63];
    end 
  end


  always @(posedge clk) begin
    if(T47) begin
      T139[0] <= io_a[62];
    end 
  end


  always @(posedge clk) begin
    if(T47) begin
      specialCodeA_PA[0] <= io_a[61];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      sign_PC <= T57;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      sign_PB <= T60;
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      sign_PA <= sign_S;
    end 
  end


  always @(posedge clk) begin
    if(N175) begin
      valid_PC <= N176;
    end 
  end


  always @(posedge clk) begin
    if(N179) begin
      cycleNum_C[2] <= N182;
    end 
  end


  always @(posedge clk) begin
    if(N179) begin
      cycleNum_C[1] <= N181;
    end 
  end


  always @(posedge clk) begin
    if(N179) begin
      cycleNum_C[0] <= N180;
    end 
  end


  always @(posedge clk) begin
    if(N185) begin
      cycleNum_B[3] <= N189;
    end 
  end


  always @(posedge clk) begin
    if(N185) begin
      cycleNum_B[2] <= N188;
    end 
  end


  always @(posedge clk) begin
    if(N185) begin
      cycleNum_B[1] <= N187;
    end 
  end


  always @(posedge clk) begin
    if(N185) begin
      cycleNum_B[0] <= N186;
    end 
  end


  always @(posedge clk) begin
    if(N192) begin
      cycleNum_A[2] <= N195;
    end 
  end


  always @(posedge clk) begin
    if(N192) begin
      cycleNum_A[1] <= N194;
    end 
  end


  always @(posedge clk) begin
    if(N192) begin
      cycleNum_A[0] <= N193;
    end 
  end


  always @(posedge clk) begin
    if(N198) begin
      valid_PA <= N199;
    end 
  end


  always @(posedge clk) begin
    if(N202) begin
      valid_PB <= N203;
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[50] <= fractB_other_PB[50];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[49] <= fractB_other_PB[49];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[48] <= fractB_other_PB[48];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[47] <= fractB_other_PB[47];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[46] <= fractB_other_PB[46];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[45] <= fractB_other_PB[45];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[44] <= fractB_other_PB[44];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[43] <= fractB_other_PB[43];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[42] <= fractB_other_PB[42];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[41] <= fractB_other_PB[41];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[40] <= fractB_other_PB[40];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[39] <= fractB_other_PB[39];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[38] <= fractB_other_PB[38];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[37] <= fractB_other_PB[37];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[36] <= fractB_other_PB[36];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[35] <= fractB_other_PB[35];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[34] <= fractB_other_PB[34];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[33] <= fractB_other_PB[33];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[32] <= fractB_other_PB[32];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[31] <= fractB_other_PB[31];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[30] <= fractB_other_PB[30];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[29] <= fractB_other_PB[29];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[28] <= fractB_other_PB[28];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[27] <= fractB_other_PB[27];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[26] <= fractB_other_PB[26];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[25] <= fractB_other_PB[25];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[24] <= fractB_other_PB[24];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[23] <= fractB_other_PB[23];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[22] <= fractB_other_PB[22];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[21] <= fractB_other_PB[21];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[20] <= fractB_other_PB[20];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[19] <= fractB_other_PB[19];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[18] <= fractB_other_PB[18];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[17] <= fractB_other_PB[17];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[16] <= fractB_other_PB[16];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[15] <= fractB_other_PB[15];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[14] <= fractB_other_PB[14];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[13] <= fractB_other_PB[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[12] <= fractB_other_PB[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[11] <= fractB_other_PB[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[10] <= fractB_other_PB[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[9] <= fractB_other_PB[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[8] <= fractB_other_PB[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[7] <= fractB_other_PB[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[6] <= fractB_other_PB[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[5] <= fractB_other_PB[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[4] <= fractB_other_PB[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[3] <= fractB_other_PB[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[2] <= fractB_other_PB[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      sigB_PC[1] <= fractB_other_PB[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T170[0] <= fractB_other_PB[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[50] <= sigB_PA_50;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[49] <= sigB_PA_49;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[48] <= sigB_PA_48;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[47] <= sigB_PA_47;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[46] <= T285[20];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[45] <= T285[19];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[44] <= T285[18];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[43] <= T285[17];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[42] <= T285[16];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[41] <= T285[15];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[40] <= T285[14];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[39] <= T285[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[38] <= T285[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[37] <= T285[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[36] <= T285[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[35] <= T285[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[34] <= T285[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[33] <= T285[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[32] <= T285[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[31] <= T285[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[30] <= T285[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[29] <= T285[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[28] <= T285[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[27] <= T285[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[26] <= T285[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[25] <= sigB_PA[25];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[24] <= sigB_PA[24];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[23] <= sigB_PA[23];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[22] <= sigB_PA[22];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[21] <= sigB_PA[21];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[20] <= sigB_PA[20];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[19] <= sigB_PA[19];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[18] <= sigB_PA[18];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[17] <= sigB_PA[17];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[16] <= sigB_PA[16];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[15] <= sigB_PA[15];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[14] <= sigB_PA[14];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[13] <= sigB_PA[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[12] <= sigB_PA[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[11] <= sigB_PA[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[10] <= sigB_PA[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[9] <= sigB_PA[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[8] <= sigB_PA[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[7] <= sigB_PA[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[6] <= sigB_PA[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[5] <= sigB_PA[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[4] <= sigB_PA[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[3] <= sigB_PA[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[2] <= sigB_PA[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[1] <= sigB_PA[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractB_other_PB[0] <= sigB_PA[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA_50 <= io_b[50];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA_49 <= io_b[49];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA_48 <= io_b[48];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA_47 <= io_b[47];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[20] <= io_b[46];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[19] <= io_b[45];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[18] <= io_b[44];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[17] <= io_b[43];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[16] <= io_b[42];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[15] <= io_b[41];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[14] <= io_b[40];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[13] <= io_b[39];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[12] <= io_b[38];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[11] <= io_b[37];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[10] <= io_b[36];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[9] <= io_b[35];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[8] <= io_b[34];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[7] <= io_b[33];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[6] <= io_b[32];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[5] <= io_b[31];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[4] <= io_b[30];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[3] <= io_b[29];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[2] <= io_b[28];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[1] <= io_b[27];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      T285[0] <= io_b[26];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[25] <= io_b[25];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[24] <= io_b[24];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[23] <= io_b[23];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[22] <= io_b[22];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[21] <= io_b[21];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[20] <= io_b[20];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[19] <= io_b[19];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[18] <= io_b[18];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[17] <= io_b[17];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[16] <= io_b[16];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[15] <= io_b[15];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[14] <= io_b[14];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[13] <= io_b[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[12] <= io_b[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[11] <= io_b[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[10] <= io_b[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[9] <= io_b[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[8] <= io_b[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[7] <= io_b[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[6] <= io_b[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[5] <= io_b[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[4] <= io_b[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[3] <= io_b[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[2] <= io_b[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[1] <= io_b[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      sigB_PA[0] <= io_b[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      sigB_PC[51] <= T180;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      fractB_51_PB <= T183;
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      sigB_PA_51 <= io_b[51];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[12] <= exp_PB[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[11] <= exp_PB[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[10] <= exp_PB[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[9] <= exp_PB[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[8] <= exp_PB[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[7] <= exp_PB[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[6] <= exp_PB[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[5] <= exp_PB[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[4] <= exp_PB[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[3] <= exp_PB[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[2] <= exp_PB[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[1] <= exp_PB[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T593[0] <= exp_PB[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      exp_PC[0] <= exp_PB[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[13] <= exp_PA[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[12] <= exp_PA[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[11] <= exp_PA[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[10] <= exp_PA[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[9] <= exp_PA[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[8] <= exp_PA[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[7] <= exp_PA[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[6] <= exp_PA[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[5] <= exp_PA[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[4] <= exp_PA[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[3] <= exp_PA[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[2] <= exp_PA[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[1] <= exp_PA[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      exp_PB[0] <= exp_PA[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[13] <= T196[13];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[12] <= T196[12];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[11] <= T196[11];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[10] <= T196[10];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[9] <= T196[9];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[8] <= T196[8];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[7] <= T196[7];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[6] <= T196[6];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[5] <= T196[5];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[4] <= T196[4];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[3] <= T196[3];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[2] <= T196[2];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[1] <= T196[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA_normalCase) begin
      exp_PA[0] <= T196[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC_normalCase) begin
      T206[53] <= fractA_0_PB;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB_normalCase) begin
      fractA_0_PB <= sigA_PA[0];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[50] <= io_a[50];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[49] <= io_a[49];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[48] <= io_a[48];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[47] <= io_a[47];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[46] <= io_a[46];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[45] <= io_a[45];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[44] <= io_a[44];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[43] <= io_a[43];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[42] <= io_a[42];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[41] <= io_a[41];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[40] <= io_a[40];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[39] <= io_a[39];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[38] <= io_a[38];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[37] <= io_a[37];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[36] <= io_a[36];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[35] <= io_a[35];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[34] <= io_a[34];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[33] <= io_a[33];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[32] <= io_a[32];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[31] <= io_a[31];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[30] <= io_a[30];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[29] <= io_a[29];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[28] <= io_a[28];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[27] <= io_a[27];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[26] <= io_a[26];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[25] <= io_a[25];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[24] <= io_a[24];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[23] <= io_a[23];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[22] <= io_a[22];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[21] <= io_a[21];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[20] <= io_a[20];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[19] <= io_a[19];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[18] <= io_a[18];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[17] <= io_a[17];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[16] <= io_a[16];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[15] <= io_a[15];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[14] <= io_a[14];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[13] <= io_a[13];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[12] <= io_a[12];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[11] <= io_a[11];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[10] <= io_a[10];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[9] <= io_a[9];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[8] <= io_a[8];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[7] <= io_a[7];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[6] <= io_a[6];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[5] <= io_a[5];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[4] <= io_a[4];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[3] <= io_a[3];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[2] <= io_a[2];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[1] <= io_a[1];
    end 
  end


  always @(posedge clk) begin
    if(T305[20]) begin
      sigA_PA[0] <= io_a[0];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      E_E_div <= E_C1_div;
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[104] <= io_mulAddResult_3[104];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[103] <= io_mulAddResult_3[103];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[102] <= io_mulAddResult_3[102];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[101] <= io_mulAddResult_3[101];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[100] <= io_mulAddResult_3[100];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[99] <= io_mulAddResult_3[99];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[98] <= io_mulAddResult_3[98];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[97] <= io_mulAddResult_3[97];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[96] <= io_mulAddResult_3[96];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[95] <= io_mulAddResult_3[95];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[94] <= io_mulAddResult_3[94];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[93] <= io_mulAddResult_3[93];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[92] <= io_mulAddResult_3[92];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[91] <= io_mulAddResult_3[91];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[90] <= io_mulAddResult_3[90];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[89] <= io_mulAddResult_3[89];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[88] <= io_mulAddResult_3[88];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[87] <= io_mulAddResult_3[87];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[86] <= io_mulAddResult_3[86];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[85] <= io_mulAddResult_3[85];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[84] <= io_mulAddResult_3[84];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[83] <= io_mulAddResult_3[83];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[82] <= io_mulAddResult_3[82];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[81] <= io_mulAddResult_3[81];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[80] <= io_mulAddResult_3[80];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[79] <= io_mulAddResult_3[79];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[78] <= io_mulAddResult_3[78];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[77] <= io_mulAddResult_3[77];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[76] <= io_mulAddResult_3[76];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[75] <= io_mulAddResult_3[75];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[74] <= io_mulAddResult_3[74];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[73] <= io_mulAddResult_3[73];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[72] <= io_mulAddResult_3[72];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[71] <= io_mulAddResult_3[71];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[70] <= io_mulAddResult_3[70];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[69] <= io_mulAddResult_3[69];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[68] <= io_mulAddResult_3[68];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[67] <= io_mulAddResult_3[67];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[66] <= io_mulAddResult_3[66];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[65] <= io_mulAddResult_3[65];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[64] <= io_mulAddResult_3[64];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[63] <= io_mulAddResult_3[63];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[62] <= io_mulAddResult_3[62];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[61] <= io_mulAddResult_3[61];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[60] <= io_mulAddResult_3[60];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[59] <= io_mulAddResult_3[59];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[58] <= io_mulAddResult_3[58];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[57] <= io_mulAddResult_3[57];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[56] <= io_mulAddResult_3[56];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[55] <= io_mulAddResult_3[55];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[54] <= io_mulAddResult_3[54];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[53] <= io_mulAddResult_3[53];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[52] <= io_mulAddResult_3[52];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[51] <= io_mulAddResult_3[51];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[50] <= io_mulAddResult_3[50];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[49] <= io_mulAddResult_3[49];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[48] <= io_mulAddResult_3[48];
    end 
  end


  always @(posedge clk) begin
    if(T221) begin
      T218[47] <= io_mulAddResult_3[47];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[103] <= io_mulAddResult_3[104];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[102] <= io_mulAddResult_3[103];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[101] <= io_mulAddResult_3[102];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[100] <= io_mulAddResult_3[101];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[99] <= io_mulAddResult_3[100];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[98] <= io_mulAddResult_3[99];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[97] <= io_mulAddResult_3[98];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[96] <= io_mulAddResult_3[97];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[95] <= io_mulAddResult_3[96];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[94] <= io_mulAddResult_3[95];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[93] <= io_mulAddResult_3[94];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[92] <= io_mulAddResult_3[93];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[91] <= io_mulAddResult_3[92];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[90] <= io_mulAddResult_3[91];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[89] <= io_mulAddResult_3[90];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[88] <= io_mulAddResult_3[89];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[87] <= io_mulAddResult_3[88];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[86] <= io_mulAddResult_3[87];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[85] <= io_mulAddResult_3[86];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[84] <= io_mulAddResult_3[85];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[83] <= io_mulAddResult_3[84];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[82] <= io_mulAddResult_3[83];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[81] <= io_mulAddResult_3[82];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[80] <= io_mulAddResult_3[81];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[79] <= io_mulAddResult_3[80];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[78] <= io_mulAddResult_3[79];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[77] <= io_mulAddResult_3[78];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[76] <= io_mulAddResult_3[77];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[75] <= io_mulAddResult_3[76];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[74] <= io_mulAddResult_3[75];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[73] <= io_mulAddResult_3[74];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[72] <= io_mulAddResult_3[73];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[71] <= io_mulAddResult_3[72];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[70] <= io_mulAddResult_3[71];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[69] <= io_mulAddResult_3[70];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[68] <= io_mulAddResult_3[69];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[67] <= io_mulAddResult_3[68];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[66] <= io_mulAddResult_3[67];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[65] <= io_mulAddResult_3[66];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[64] <= io_mulAddResult_3[65];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[63] <= io_mulAddResult_3[64];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[62] <= io_mulAddResult_3[63];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[61] <= io_mulAddResult_3[62];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[60] <= io_mulAddResult_3[61];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[59] <= io_mulAddResult_3[60];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[58] <= io_mulAddResult_3[59];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[57] <= io_mulAddResult_3[58];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[56] <= io_mulAddResult_3[57];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[55] <= io_mulAddResult_3[56];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[54] <= io_mulAddResult_3[55];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[53] <= io_mulAddResult_3[54];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[52] <= io_mulAddResult_3[53];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[51] <= io_mulAddResult_3[52];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[50] <= io_mulAddResult_3[51];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[49] <= io_mulAddResult_3[50];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[48] <= io_mulAddResult_3[49];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[47] <= io_mulAddResult_3[48];
    end 
  end


  always @(posedge clk) begin
    if(N493) begin
      T230[46] <= io_mulAddResult_3[47];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      sqrSigma1_C[32] <= io_mulAddResult_3[79];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      sqrSigma1_C[31] <= io_mulAddResult_3[78];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[29] <= io_mulAddResult_3[77];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[28] <= io_mulAddResult_3[76];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[27] <= io_mulAddResult_3[75];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[26] <= io_mulAddResult_3[74];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[25] <= io_mulAddResult_3[73];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[24] <= io_mulAddResult_3[72];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[23] <= io_mulAddResult_3[71];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[22] <= io_mulAddResult_3[70];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[21] <= io_mulAddResult_3[69];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[20] <= io_mulAddResult_3[68];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[19] <= io_mulAddResult_3[67];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[18] <= io_mulAddResult_3[66];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[17] <= io_mulAddResult_3[65];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[16] <= io_mulAddResult_3[64];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[15] <= io_mulAddResult_3[63];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[14] <= io_mulAddResult_3[62];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[13] <= io_mulAddResult_3[61];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[12] <= io_mulAddResult_3[60];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[11] <= io_mulAddResult_3[59];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[10] <= io_mulAddResult_3[58];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[9] <= io_mulAddResult_3[57];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[8] <= io_mulAddResult_3[56];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[7] <= io_mulAddResult_3[55];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[6] <= io_mulAddResult_3[54];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[5] <= io_mulAddResult_3[53];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[4] <= io_mulAddResult_3[52];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[3] <= io_mulAddResult_3[51];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[2] <= io_mulAddResult_3[50];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[1] <= io_mulAddResult_3[49];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      T241[0] <= io_mulAddResult_3[48];
    end 
  end


  always @(posedge clk) begin
    if(N489) begin
      sqrSigma1_C_0 <= io_mulAddResult_3[47];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[52] <= ER1_A1_sqrt[16];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[51] <= ER1_A1_sqrt[15];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[50] <= ER1_A1_sqrt[14];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[49] <= ER1_A1_sqrt[13];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[48] <= ER1_A1_sqrt[12];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[47] <= ER1_A1_sqrt[11];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[46] <= ER1_A1_sqrt[10];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[45] <= ER1_A1_sqrt[9];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[44] <= ER1_A1_sqrt[8];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[43] <= ER1_A1_sqrt[7];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[42] <= ER1_A1_sqrt[6];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[41] <= ER1_A1_sqrt[5];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[40] <= ER1_A1_sqrt[4];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[39] <= ER1_A1_sqrt[3];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[38] <= ER1_A1_sqrt[2];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[37] <= ER1_A1_sqrt[1];
    end 
  end


  always @(posedge clk) begin
    if(cyc_A1_sqrt) begin
      T248[36] <= ER1_A1_sqrt[0];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[23] <= T258[8];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[22] <= T258[7];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[21] <= T258[6];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[20] <= T258[5];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[19] <= T258[4];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[18] <= T258[3];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[17] <= T258[2];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[16] <= T258[1];
    end 
  end


  always @(posedge clk) begin
    if(T269) begin
      T256[15] <= T258[0];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[20] <= T277[20];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[19] <= T277[19];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[18] <= T277[18];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[17] <= T277[17];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[16] <= T277[16];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[15] <= T277[15];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[14] <= T277[14];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[13] <= T277[13];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[12] <= T277[12];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[11] <= T277[11];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[10] <= T277[10];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[9] <= T277[9];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[8] <= T277[8];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[7] <= T277[7];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[6] <= T277[6];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[5] <= T277[5];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[4] <= T277[4];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[3] <= T277[3];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[2] <= T277[2];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[1] <= T277[1];
    end 
  end


  always @(posedge clk) begin
    if(T280) begin
      partNegSigma0_A[0] <= T277[0];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[9] <= T292[9];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[8] <= T292[8];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[7] <= T292[7];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[6] <= T292[6];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[5] <= T292[5];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[4] <= T292[4];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[3] <= T292[3];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[2] <= T292[2];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[1] <= T292[1];
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      T908[0] <= T292[0];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[8] <= T390[8];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[7] <= T390[7];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[6] <= T390[6];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[5] <= T390[5];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[4] <= T390[4];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[3] <= T390[3];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[2] <= T390[2];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[1] <= T390[1];
    end 
  end


  always @(posedge clk) begin
    if(T403) begin
      nextMulAdd9B_A[0] <= T390[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[8] <= T917[8];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[7] <= T917[7];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[6] <= T917[6];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[5] <= T917[5];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[4] <= T917[4];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[3] <= T917[3];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[2] <= T917[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[1] <= T917[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T918[0] <= T917[0];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[50] <= io_mulAddResult_3[103];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[49] <= io_mulAddResult_3[102];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[48] <= io_mulAddResult_3[101];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[47] <= io_mulAddResult_3[100];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[46] <= io_mulAddResult_3[99];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[45] <= io_mulAddResult_3[98];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[44] <= io_mulAddResult_3[97];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[43] <= io_mulAddResult_3[96];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[42] <= io_mulAddResult_3[95];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[41] <= io_mulAddResult_3[94];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[40] <= io_mulAddResult_3[93];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[39] <= io_mulAddResult_3[92];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[38] <= io_mulAddResult_3[91];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[37] <= io_mulAddResult_3[90];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[36] <= io_mulAddResult_3[89];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[35] <= io_mulAddResult_3[88];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[34] <= io_mulAddResult_3[87];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[33] <= io_mulAddResult_3[86];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[32] <= io_mulAddResult_3[85];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[31] <= io_mulAddResult_3[84];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[30] <= io_mulAddResult_3[83];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[29] <= io_mulAddResult_3[82];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[28] <= io_mulAddResult_3[81];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[27] <= io_mulAddResult_3[80];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[26] <= io_mulAddResult_3[79];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[25] <= io_mulAddResult_3[78];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[24] <= io_mulAddResult_3[77];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[23] <= io_mulAddResult_3[76];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[22] <= io_mulAddResult_3[75];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[21] <= io_mulAddResult_3[74];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[20] <= io_mulAddResult_3[73];
    end 
  end


  always @(posedge clk) begin
    if(N294) begin
      T472[19] <= io_mulAddResult_3[72];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[45] <= io_mulAddResult_3[103];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[44] <= io_mulAddResult_3[102];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[43] <= io_mulAddResult_3[101];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[42] <= io_mulAddResult_3[100];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[41] <= io_mulAddResult_3[99];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[40] <= io_mulAddResult_3[98];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[39] <= io_mulAddResult_3[97];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[38] <= io_mulAddResult_3[96];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[37] <= io_mulAddResult_3[95];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[36] <= io_mulAddResult_3[94];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[35] <= io_mulAddResult_3[93];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[34] <= io_mulAddResult_3[92];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[33] <= io_mulAddResult_3[91];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[32] <= io_mulAddResult_3[90];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[31] <= io_mulAddResult_3[89];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[30] <= io_mulAddResult_3[88];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[29] <= io_mulAddResult_3[87];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[28] <= io_mulAddResult_3[86];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[27] <= io_mulAddResult_3[85];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[26] <= io_mulAddResult_3[84];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[25] <= io_mulAddResult_3[83];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[24] <= io_mulAddResult_3[82];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[23] <= io_mulAddResult_3[81];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[22] <= io_mulAddResult_3[80];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[21] <= io_mulAddResult_3[79];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[20] <= io_mulAddResult_3[78];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[19] <= io_mulAddResult_3[77];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[18] <= io_mulAddResult_3[76];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[17] <= io_mulAddResult_3[75];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[16] <= io_mulAddResult_3[74];
    end 
  end


  always @(posedge clk) begin
    if(cyc_C5_sqrt) begin
      T491[15] <= io_mulAddResult_3[73];
    end 
  end


  always @(posedge clk) begin
    if(T47) begin
      sigA_PA[51] <= io_a[51];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[52] <= sigT_C1[53];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[51] <= sigT_C1[52];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[50] <= sigT_C1[51];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[49] <= sigT_C1[50];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[48] <= sigT_C1[49];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[47] <= sigT_C1[48];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[46] <= sigT_C1[47];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[45] <= sigT_C1[46];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[44] <= sigT_C1[45];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[43] <= sigT_C1[44];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[42] <= sigT_C1[43];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[41] <= sigT_C1[42];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[40] <= sigT_C1[41];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[39] <= sigT_C1[40];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[38] <= sigT_C1[39];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[37] <= sigT_C1[38];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[36] <= sigT_C1[37];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[35] <= sigT_C1[36];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[34] <= sigT_C1[35];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[33] <= sigT_C1[34];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[32] <= sigT_C1[33];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[31] <= sigT_C1[32];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[30] <= sigT_C1[31];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[29] <= sigT_C1[30];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[28] <= sigT_C1[29];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[27] <= sigT_C1[28];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[26] <= sigT_C1[27];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[25] <= sigT_C1[26];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[24] <= sigT_C1[25];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[23] <= sigT_C1[24];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[22] <= sigT_C1[23];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[21] <= sigT_C1[22];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[20] <= sigT_C1[21];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[19] <= sigT_C1[20];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[18] <= sigT_C1[19];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[17] <= sigT_C1[18];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[16] <= sigT_C1[17];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[15] <= sigT_C1[16];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[14] <= sigT_C1[15];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[13] <= sigT_C1[14];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[12] <= sigT_C1[13];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[11] <= sigT_C1[12];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[10] <= sigT_C1[11];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[9] <= sigT_C1[10];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[8] <= sigT_C1[9];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[7] <= sigT_C1[8];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[6] <= sigT_C1[7];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[5] <= sigT_C1[6];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[4] <= sigT_C1[5];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[3] <= sigT_C1[4];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[2] <= sigT_C1[3];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[1] <= sigT_C1[2];
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T727[0] <= sigT_C1[1];
    end 
  end


  always @(posedge clk) begin
    if(N272) begin
      isZeroRemT_E <= T680;
    end 
  end


  always @(posedge clk) begin
    if(N272) begin
      isNegRemT_E <= T693;
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      roundingMode_PC[1] <= T720[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      roundingMode_PC[0] <= T720[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      roundingMode_PB[1] <= T722[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      roundingMode_PB[0] <= T722[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      roundingMode_PA[1] <= io_roundingMode[1];
    end 
  end


  always @(posedge clk) begin
    if(entering_PA) begin
      roundingMode_PA[0] <= io_roundingMode[0];
    end 
  end


  always @(posedge clk) begin
    if(entering_PC) begin
      fractA_51_PC <= T803;
    end 
  end


  always @(posedge clk) begin
    if(entering_PB) begin
      fractA_51_PB <= T806;
    end 
  end

  assign N213 = io_mulAddResult_3[52] | io_mulAddResult_3[53];
  assign N214 = io_mulAddResult_3[51] | N213;
  assign N215 = io_mulAddResult_3[50] | N214;
  assign N216 = io_mulAddResult_3[49] | N215;
  assign N217 = io_mulAddResult_3[48] | N216;
  assign N218 = io_mulAddResult_3[47] | N217;
  assign N219 = io_mulAddResult_3[46] | N218;
  assign N220 = io_mulAddResult_3[45] | N219;
  assign N221 = io_mulAddResult_3[44] | N220;
  assign N222 = io_mulAddResult_3[43] | N221;
  assign N223 = io_mulAddResult_3[42] | N222;
  assign N224 = io_mulAddResult_3[41] | N223;
  assign N225 = io_mulAddResult_3[40] | N224;
  assign N226 = io_mulAddResult_3[39] | N225;
  assign N227 = io_mulAddResult_3[38] | N226;
  assign N228 = io_mulAddResult_3[37] | N227;
  assign N229 = io_mulAddResult_3[36] | N228;
  assign N230 = io_mulAddResult_3[35] | N229;
  assign N231 = io_mulAddResult_3[34] | N230;
  assign N232 = io_mulAddResult_3[33] | N231;
  assign N233 = io_mulAddResult_3[32] | N232;
  assign N234 = io_mulAddResult_3[31] | N233;
  assign N235 = io_mulAddResult_3[30] | N234;
  assign N236 = io_mulAddResult_3[29] | N235;
  assign N237 = io_mulAddResult_3[28] | N236;
  assign N238 = io_mulAddResult_3[27] | N237;
  assign N239 = io_mulAddResult_3[26] | N238;
  assign N240 = io_mulAddResult_3[25] | N239;
  assign N241 = io_mulAddResult_3[24] | N240;
  assign N242 = io_mulAddResult_3[23] | N241;
  assign N243 = io_mulAddResult_3[22] | N242;
  assign N244 = io_mulAddResult_3[21] | N243;
  assign N245 = io_mulAddResult_3[20] | N244;
  assign N246 = io_mulAddResult_3[19] | N245;
  assign N247 = io_mulAddResult_3[18] | N246;
  assign N248 = io_mulAddResult_3[17] | N247;
  assign N249 = io_mulAddResult_3[16] | N248;
  assign N250 = io_mulAddResult_3[15] | N249;
  assign N251 = io_mulAddResult_3[14] | N250;
  assign N252 = io_mulAddResult_3[13] | N251;
  assign N253 = io_mulAddResult_3[12] | N252;
  assign N254 = io_mulAddResult_3[11] | N253;
  assign N255 = io_mulAddResult_3[10] | N254;
  assign N256 = io_mulAddResult_3[9] | N255;
  assign N257 = io_mulAddResult_3[8] | N256;
  assign N258 = io_mulAddResult_3[7] | N257;
  assign N259 = io_mulAddResult_3[6] | N258;
  assign N260 = io_mulAddResult_3[5] | N259;
  assign N261 = io_mulAddResult_3[4] | N260;
  assign N262 = io_mulAddResult_3[3] | N261;
  assign N263 = io_mulAddResult_3[2] | N262;
  assign N264 = io_mulAddResult_3[1] | N263;
  assign N265 = io_mulAddResult_3[0] | N264;
  assign N266 = ~N265;
  assign N267 = io_mulAddResult_3[54] | io_mulAddResult_3[55];
  assign N268 = ~N267;
  assign N269 = ~cycleNum_E[1];
  assign N270 = N269 | cycleNum_E[2];
  assign N271 = cycleNum_E[0] | N270;
  assign N272 = ~N271;
  assign N273 = cycleNum_E[1] | cycleNum_E[2];
  assign N274 = cycleNum_E[0] | N273;
  assign N275 = cycleNum_C[1] | cycleNum_C[2];
  assign N276 = cycleNum_C[0] | N275;
  assign N277 = cycleNum_B[2] | cycleNum_B[3];
  assign N278 = cycleNum_B[1] | N277;
  assign N279 = cycleNum_B[0] | N278;
  assign N280 = cycleNum_A[1] | cycleNum_A[2];
  assign N281 = cycleNum_A[0] | N280;
  assign N282 = ~cycleNum_C[1];
  assign N283 = N282 | cycleNum_C[2];
  assign N284 = cycleNum_C[0] | N283;
  assign N285 = ~N284;
  assign N286 = ~cycleNum_E[0];
  assign N287 = N269 | cycleNum_E[2];
  assign N288 = N286 | N287;
  assign N289 = ~N288;
  assign N290 = ~cycleNum_B[3];
  assign N291 = cycleNum_B[2] | N290;
  assign N292 = cycleNum_B[1] | N291;
  assign N293 = cycleNum_B[0] | N292;
  assign N294 = ~N293;
  assign N295 = ~cycleNum_B[1];
  assign N296 = cycleNum_B[2] | N290;
  assign N297 = N295 | N296;
  assign N298 = cycleNum_B[0] | N297;
  assign N299 = ~N298;
  assign N300 = ~cycleNum_B[0];
  assign N301 = cycleNum_B[2] | N290;
  assign N302 = cycleNum_B[1] | N301;
  assign N303 = N300 | N302;
  assign N304 = ~N303;
  assign N305 = ~cycleNum_C[2];
  assign N306 = N282 | N305;
  assign N307 = cycleNum_C[0] | N306;
  assign N308 = ~N307;
  assign N309 = ~cycleNum_C[0];
  assign N310 = cycleNum_C[1] | cycleNum_C[2];
  assign N311 = N309 | N310;
  assign N312 = ~N311;
  assign N313 = ~cycleNum_A[0];
  assign N314 = cycleNum_A[1] | cycleNum_A[2];
  assign N315 = N313 | N314;
  assign N316 = ~N315;
  assign N317 = ~cycleNum_A[1];
  assign N318 = N317 | cycleNum_A[2];
  assign N319 = cycleNum_A[0] | N318;
  assign N320 = ~N319;
  assign N321 = ~cycleNum_A[2];
  assign N322 = cycleNum_A[1] | N321;
  assign N323 = N313 | N322;
  assign N324 = ~N323;
  assign N325 = cycleNum_A[1] | N321;
  assign N326 = cycleNum_A[0] | N325;
  assign N327 = ~N326;
  assign N328 = N317 | cycleNum_A[2];
  assign N329 = N313 | N328;
  assign N330 = ~N329;
  assign N331 = io_b[50] & io_b[51];
  assign N332 = io_b[49] & N331;
  assign N333 = ~io_b[51];
  assign N334 = ~io_b[50];
  assign N335 = N334 | N333;
  assign N336 = io_b[49] | N335;
  assign N337 = ~N336;
  assign N338 = ~io_b[49];
  assign N339 = io_b[50] | N333;
  assign N340 = N338 | N339;
  assign N341 = ~N340;
  assign N342 = io_b[49] | N339;
  assign N343 = ~N342;
  assign N344 = N334 | io_b[51];
  assign N345 = N338 | N344;
  assign N346 = ~N345;
  assign N347 = N317 | N321;
  assign N348 = cycleNum_A[0] | N347;
  assign N349 = ~N348;
  assign N350 = io_b[49] | N344;
  assign N351 = ~N350;
  assign N352 = io_b[50] | io_b[51];
  assign N353 = io_b[49] | N352;
  assign N354 = ~N353;
  assign N355 = N338 | N352;
  assign N356 = ~N355;
  assign N357 = T581[51] | T581[52];
  assign N358 = T581[50] | N357;
  assign N359 = T581[49] | N358;
  assign N360 = T581[48] | N359;
  assign N361 = T581[47] | N360;
  assign N362 = T581[46] | N361;
  assign N363 = T581[45] | N362;
  assign N364 = T581[44] | N363;
  assign N365 = T581[43] | N364;
  assign N366 = T581[42] | N365;
  assign N367 = T581[41] | N366;
  assign N368 = T581[40] | N367;
  assign N369 = T581[39] | N368;
  assign N370 = T581[38] | N369;
  assign N371 = T581[37] | N370;
  assign N372 = T581[36] | N371;
  assign N373 = T581[35] | N372;
  assign N374 = T581[34] | N373;
  assign N375 = T581[33] | N374;
  assign N376 = T581[32] | N375;
  assign N377 = T581[31] | N376;
  assign N378 = T581[30] | N377;
  assign N379 = T581[29] | N378;
  assign N380 = T581[28] | N379;
  assign N381 = T581[27] | N380;
  assign N382 = T581[26] | N381;
  assign N383 = T581[25] | N382;
  assign N384 = T581[24] | N383;
  assign N385 = T581[23] | N384;
  assign N386 = T581[22] | N385;
  assign N387 = T581[21] | N386;
  assign N388 = T581[20] | N387;
  assign N389 = T581[19] | N388;
  assign N390 = T581[18] | N389;
  assign N391 = T581[17] | N390;
  assign N392 = T581[16] | N391;
  assign N393 = T581[15] | N392;
  assign N394 = T581[14] | N393;
  assign N395 = T581[13] | N394;
  assign N396 = T581[12] | N395;
  assign N397 = T581[11] | N396;
  assign N398 = T581[10] | N397;
  assign N399 = T581[9] | N398;
  assign N400 = T581[8] | N399;
  assign N401 = T581[7] | N400;
  assign N402 = T581[6] | N401;
  assign N403 = T581[5] | N402;
  assign N404 = T581[4] | N403;
  assign N405 = T581[3] | N404;
  assign N406 = T581[2] | N405;
  assign N407 = T581[1] | N406;
  assign N408 = T581[0] | N407;
  assign N409 = ~N408;
  assign N410 = roundingMode_PC[0] | roundingMode_PC[1];
  assign N411 = ~N410;
  assign N412 = T700[51] | T700[52];
  assign N413 = T700[50] | N412;
  assign N414 = T700[49] | N413;
  assign N415 = T700[48] | N414;
  assign N416 = T700[47] | N415;
  assign N417 = T700[46] | N416;
  assign N418 = T700[45] | N417;
  assign N419 = T700[44] | N418;
  assign N420 = T700[43] | N419;
  assign N421 = T700[42] | N420;
  assign N422 = T700[41] | N421;
  assign N423 = T700[40] | N422;
  assign N424 = T700[39] | N423;
  assign N425 = T700[38] | N424;
  assign N426 = T700[37] | N425;
  assign N427 = T700[36] | N426;
  assign N428 = T700[35] | N427;
  assign N429 = T700[34] | N428;
  assign N430 = T700[33] | N429;
  assign N431 = T700[32] | N430;
  assign N432 = T700[31] | N431;
  assign N433 = T700[30] | N432;
  assign N434 = T700[29] | N433;
  assign N435 = T700[28] | N434;
  assign N436 = T700[27] | N435;
  assign N437 = T700[26] | N436;
  assign N438 = T700[25] | N437;
  assign N439 = T700[24] | N438;
  assign N440 = T700[23] | N439;
  assign N441 = T700[22] | N440;
  assign N442 = T700[21] | N441;
  assign N443 = T700[20] | N442;
  assign N444 = T700[19] | N443;
  assign N445 = T700[18] | N444;
  assign N446 = T700[17] | N445;
  assign N447 = T700[16] | N446;
  assign N448 = T700[15] | N447;
  assign N449 = T700[14] | N448;
  assign N450 = T700[13] | N449;
  assign N451 = T700[12] | N450;
  assign N452 = T700[11] | N451;
  assign N453 = T700[10] | N452;
  assign N454 = T700[9] | N453;
  assign N455 = T700[8] | N454;
  assign N456 = T700[7] | N455;
  assign N457 = T700[6] | N456;
  assign N458 = T700[5] | N457;
  assign N459 = T700[4] | N458;
  assign N460 = T700[3] | N459;
  assign N461 = T700[2] | N460;
  assign N462 = T700[1] | N461;
  assign N463 = T700[0] | N462;
  assign N464 = io_b[62] | io_b[63];
  assign N465 = io_b[61] | N464;
  assign N466 = ~N465;
  assign N467 = ~roundingMode_PC[1];
  assign N468 = roundingMode_PC[0] | N467;
  assign N469 = ~N468;
  assign N470 = roundingMode_PC[0] & roundingMode_PC[1];
  assign N471 = io_a[62] | io_a[63];
  assign N472 = io_a[61] | N471;
  assign N473 = ~N472;
  assign N474 = cycleNum_C[1] | N305;
  assign N475 = cycleNum_C[0] | N474;
  assign N476 = ~N475;
  assign N477 = io_a[62] & io_a[63];
  assign N478 = io_b[62] & io_b[63];
  assign N479 = cycleNum_C[1] | N305;
  assign N480 = N309 | N479;
  assign N481 = ~N480;
  assign N482 = cycleNum_B[2] | cycleNum_B[3];
  assign N483 = N295 | N482;
  assign N484 = cycleNum_B[0] | N483;
  assign N485 = ~N484;
  assign N486 = cycleNum_B[2] | cycleNum_B[3];
  assign N487 = cycleNum_B[1] | N486;
  assign N488 = N300 | N487;
  assign N489 = ~N488;
  assign N490 = cycleNum_B[2] | cycleNum_B[3];
  assign N491 = N295 | N490;
  assign N492 = N300 | N491;
  assign N493 = ~N492;
  assign { SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, SV2V_UNCONNECTED_16, SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, SV2V_UNCONNECTED_32, SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, SV2V_UNCONNECTED_49, SV2V_UNCONNECTED_50, SV2V_UNCONNECTED_51, SV2V_UNCONNECTED_52, SV2V_UNCONNECTED_53, SV2V_UNCONNECTED_54, SV2V_UNCONNECTED_55, SV2V_UNCONNECTED_56, SV2V_UNCONNECTED_57, SV2V_UNCONNECTED_58, SV2V_UNCONNECTED_59, SV2V_UNCONNECTED_60, SV2V_UNCONNECTED_61, SV2V_UNCONNECTED_62, SV2V_UNCONNECTED_63, SV2V_UNCONNECTED_64, SV2V_UNCONNECTED_65, SV2V_UNCONNECTED_66, SV2V_UNCONNECTED_67, SV2V_UNCONNECTED_68, SV2V_UNCONNECTED_69, SV2V_UNCONNECTED_70, SV2V_UNCONNECTED_71, SV2V_UNCONNECTED_72, SV2V_UNCONNECTED_73, SV2V_UNCONNECTED_74, SV2V_UNCONNECTED_75, SV2V_UNCONNECTED_76, SV2V_UNCONNECTED_77, SV2V_UNCONNECTED_78, SV2V_UNCONNECTED_79, SV2V_UNCONNECTED_80, SV2V_UNCONNECTED_81, SV2V_UNCONNECTED_82, SV2V_UNCONNECTED_83, SV2V_UNCONNECTED_84, SV2V_UNCONNECTED_85, SV2V_UNCONNECTED_86, SV2V_UNCONNECTED_87, SV2V_UNCONNECTED_88, SV2V_UNCONNECTED_89, SV2V_UNCONNECTED_90, SV2V_UNCONNECTED_91, SV2V_UNCONNECTED_92, SV2V_UNCONNECTED_93, SV2V_UNCONNECTED_94, SV2V_UNCONNECTED_95, SV2V_UNCONNECTED_96, SV2V_UNCONNECTED_97, SV2V_UNCONNECTED_98, SV2V_UNCONNECTED_99, SV2V_UNCONNECTED_100, SV2V_UNCONNECTED_101, SV2V_UNCONNECTED_102, SV2V_UNCONNECTED_103, SV2V_UNCONNECTED_104, SV2V_UNCONNECTED_105, SV2V_UNCONNECTED_106, SV2V_UNCONNECTED_107, SV2V_UNCONNECTED_108, SV2V_UNCONNECTED_109, SV2V_UNCONNECTED_110, SV2V_UNCONNECTED_111, SV2V_UNCONNECTED_112, SV2V_UNCONNECTED_113, SV2V_UNCONNECTED_114, SV2V_UNCONNECTED_115, SV2V_UNCONNECTED_116, SV2V_UNCONNECTED_117, SV2V_UNCONNECTED_118, SV2V_UNCONNECTED_119, SV2V_UNCONNECTED_120, SV2V_UNCONNECTED_121, SV2V_UNCONNECTED_122, SV2V_UNCONNECTED_123, SV2V_UNCONNECTED_124, SV2V_UNCONNECTED_125, SV2V_UNCONNECTED_126, SV2V_UNCONNECTED_127, SV2V_UNCONNECTED_128, SV2V_UNCONNECTED_129, SV2V_UNCONNECTED_130, SV2V_UNCONNECTED_131, SV2V_UNCONNECTED_132, SV2V_UNCONNECTED_133, SV2V_UNCONNECTED_134, SV2V_UNCONNECTED_135, SV2V_UNCONNECTED_136, SV2V_UNCONNECTED_137, SV2V_UNCONNECTED_138, SV2V_UNCONNECTED_139, SV2V_UNCONNECTED_140, SV2V_UNCONNECTED_141, SV2V_UNCONNECTED_142, SV2V_UNCONNECTED_143, SV2V_UNCONNECTED_144, SV2V_UNCONNECTED_145, SV2V_UNCONNECTED_146, SV2V_UNCONNECTED_147, SV2V_UNCONNECTED_148, SV2V_UNCONNECTED_149, SV2V_UNCONNECTED_150, SV2V_UNCONNECTED_151, SV2V_UNCONNECTED_152, SV2V_UNCONNECTED_153, SV2V_UNCONNECTED_154, SV2V_UNCONNECTED_155, SV2V_UNCONNECTED_156, SV2V_UNCONNECTED_157, SV2V_UNCONNECTED_158, SV2V_UNCONNECTED_159, SV2V_UNCONNECTED_160, SV2V_UNCONNECTED_161, SV2V_UNCONNECTED_162, SV2V_UNCONNECTED_163, SV2V_UNCONNECTED_164, SV2V_UNCONNECTED_165, SV2V_UNCONNECTED_166, SV2V_UNCONNECTED_167, SV2V_UNCONNECTED_168, SV2V_UNCONNECTED_169, SV2V_UNCONNECTED_170, SV2V_UNCONNECTED_171, SV2V_UNCONNECTED_172, SV2V_UNCONNECTED_173, SV2V_UNCONNECTED_174, SV2V_UNCONNECTED_175, SV2V_UNCONNECTED_176, SV2V_UNCONNECTED_177, SV2V_UNCONNECTED_178, SV2V_UNCONNECTED_179, SV2V_UNCONNECTED_180, SV2V_UNCONNECTED_181, SV2V_UNCONNECTED_182, SV2V_UNCONNECTED_183, SV2V_UNCONNECTED_184, SV2V_UNCONNECTED_185, SV2V_UNCONNECTED_186, SV2V_UNCONNECTED_187, SV2V_UNCONNECTED_188, SV2V_UNCONNECTED_189, SV2V_UNCONNECTED_190, SV2V_UNCONNECTED_191, SV2V_UNCONNECTED_192, SV2V_UNCONNECTED_193, SV2V_UNCONNECTED_194, SV2V_UNCONNECTED_195, SV2V_UNCONNECTED_196, SV2V_UNCONNECTED_197, SV2V_UNCONNECTED_198, SV2V_UNCONNECTED_199, SV2V_UNCONNECTED_200, SV2V_UNCONNECTED_201, SV2V_UNCONNECTED_202, SV2V_UNCONNECTED_203, SV2V_UNCONNECTED_204, SV2V_UNCONNECTED_205, SV2V_UNCONNECTED_206, SV2V_UNCONNECTED_207, SV2V_UNCONNECTED_208, SV2V_UNCONNECTED_209, SV2V_UNCONNECTED_210, SV2V_UNCONNECTED_211, SV2V_UNCONNECTED_212, SV2V_UNCONNECTED_213, SV2V_UNCONNECTED_214, SV2V_UNCONNECTED_215, SV2V_UNCONNECTED_216, SV2V_UNCONNECTED_217, SV2V_UNCONNECTED_218, SV2V_UNCONNECTED_219, SV2V_UNCONNECTED_220, SV2V_UNCONNECTED_221, SV2V_UNCONNECTED_222, SV2V_UNCONNECTED_223, SV2V_UNCONNECTED_224, SV2V_UNCONNECTED_225, SV2V_UNCONNECTED_226, SV2V_UNCONNECTED_227, SV2V_UNCONNECTED_228, SV2V_UNCONNECTED_229, SV2V_UNCONNECTED_230, SV2V_UNCONNECTED_231, SV2V_UNCONNECTED_232, SV2V_UNCONNECTED_233, SV2V_UNCONNECTED_234, SV2V_UNCONNECTED_235, SV2V_UNCONNECTED_236, SV2V_UNCONNECTED_237, SV2V_UNCONNECTED_238, SV2V_UNCONNECTED_239, SV2V_UNCONNECTED_240, SV2V_UNCONNECTED_241, SV2V_UNCONNECTED_242, SV2V_UNCONNECTED_243, SV2V_UNCONNECTED_244, SV2V_UNCONNECTED_245, SV2V_UNCONNECTED_246, SV2V_UNCONNECTED_247, SV2V_UNCONNECTED_248, SV2V_UNCONNECTED_249, SV2V_UNCONNECTED_250, SV2V_UNCONNECTED_251, SV2V_UNCONNECTED_252, SV2V_UNCONNECTED_253, SV2V_UNCONNECTED_254, SV2V_UNCONNECTED_255, SV2V_UNCONNECTED_256, SV2V_UNCONNECTED_257, SV2V_UNCONNECTED_258, SV2V_UNCONNECTED_259, SV2V_UNCONNECTED_260, SV2V_UNCONNECTED_261, SV2V_UNCONNECTED_262, SV2V_UNCONNECTED_263, SV2V_UNCONNECTED_264, SV2V_UNCONNECTED_265, SV2V_UNCONNECTED_266, SV2V_UNCONNECTED_267, SV2V_UNCONNECTED_268, SV2V_UNCONNECTED_269, SV2V_UNCONNECTED_270, SV2V_UNCONNECTED_271, SV2V_UNCONNECTED_272, SV2V_UNCONNECTED_273, SV2V_UNCONNECTED_274, SV2V_UNCONNECTED_275, SV2V_UNCONNECTED_276, SV2V_UNCONNECTED_277, SV2V_UNCONNECTED_278, SV2V_UNCONNECTED_279, SV2V_UNCONNECTED_280, SV2V_UNCONNECTED_281, SV2V_UNCONNECTED_282, SV2V_UNCONNECTED_283, SV2V_UNCONNECTED_284, SV2V_UNCONNECTED_285, SV2V_UNCONNECTED_286, SV2V_UNCONNECTED_287, SV2V_UNCONNECTED_288, SV2V_UNCONNECTED_289, SV2V_UNCONNECTED_290, SV2V_UNCONNECTED_291, SV2V_UNCONNECTED_292, SV2V_UNCONNECTED_293, SV2V_UNCONNECTED_294, SV2V_UNCONNECTED_295, SV2V_UNCONNECTED_296, SV2V_UNCONNECTED_297, SV2V_UNCONNECTED_298, SV2V_UNCONNECTED_299, SV2V_UNCONNECTED_300, SV2V_UNCONNECTED_301, SV2V_UNCONNECTED_302, SV2V_UNCONNECTED_303, SV2V_UNCONNECTED_304, SV2V_UNCONNECTED_305, SV2V_UNCONNECTED_306, SV2V_UNCONNECTED_307, SV2V_UNCONNECTED_308, SV2V_UNCONNECTED_309, SV2V_UNCONNECTED_310, SV2V_UNCONNECTED_311, SV2V_UNCONNECTED_312, SV2V_UNCONNECTED_313, SV2V_UNCONNECTED_314, SV2V_UNCONNECTED_315, SV2V_UNCONNECTED_316, SV2V_UNCONNECTED_317, SV2V_UNCONNECTED_318, SV2V_UNCONNECTED_319, SV2V_UNCONNECTED_320, SV2V_UNCONNECTED_321, SV2V_UNCONNECTED_322, SV2V_UNCONNECTED_323, SV2V_UNCONNECTED_324, SV2V_UNCONNECTED_325, SV2V_UNCONNECTED_326, SV2V_UNCONNECTED_327, SV2V_UNCONNECTED_328, SV2V_UNCONNECTED_329, SV2V_UNCONNECTED_330, SV2V_UNCONNECTED_331, SV2V_UNCONNECTED_332, SV2V_UNCONNECTED_333, SV2V_UNCONNECTED_334, SV2V_UNCONNECTED_335, SV2V_UNCONNECTED_336, SV2V_UNCONNECTED_337, SV2V_UNCONNECTED_338, SV2V_UNCONNECTED_339, SV2V_UNCONNECTED_340, SV2V_UNCONNECTED_341, SV2V_UNCONNECTED_342, SV2V_UNCONNECTED_343, SV2V_UNCONNECTED_344, SV2V_UNCONNECTED_345, SV2V_UNCONNECTED_346, SV2V_UNCONNECTED_347, SV2V_UNCONNECTED_348, SV2V_UNCONNECTED_349, SV2V_UNCONNECTED_350, SV2V_UNCONNECTED_351, SV2V_UNCONNECTED_352, SV2V_UNCONNECTED_353, SV2V_UNCONNECTED_354, SV2V_UNCONNECTED_355, SV2V_UNCONNECTED_356, SV2V_UNCONNECTED_357, SV2V_UNCONNECTED_358, SV2V_UNCONNECTED_359, SV2V_UNCONNECTED_360, SV2V_UNCONNECTED_361, SV2V_UNCONNECTED_362, SV2V_UNCONNECTED_363, SV2V_UNCONNECTED_364, SV2V_UNCONNECTED_365, SV2V_UNCONNECTED_366, SV2V_UNCONNECTED_367, SV2V_UNCONNECTED_368, SV2V_UNCONNECTED_369, SV2V_UNCONNECTED_370, SV2V_UNCONNECTED_371, SV2V_UNCONNECTED_372, SV2V_UNCONNECTED_373, SV2V_UNCONNECTED_374, SV2V_UNCONNECTED_375, SV2V_UNCONNECTED_376, SV2V_UNCONNECTED_377, SV2V_UNCONNECTED_378, SV2V_UNCONNECTED_379, SV2V_UNCONNECTED_380, SV2V_UNCONNECTED_381, SV2V_UNCONNECTED_382, SV2V_UNCONNECTED_383, SV2V_UNCONNECTED_384, SV2V_UNCONNECTED_385, SV2V_UNCONNECTED_386, SV2V_UNCONNECTED_387, SV2V_UNCONNECTED_388, SV2V_UNCONNECTED_389, SV2V_UNCONNECTED_390, SV2V_UNCONNECTED_391, SV2V_UNCONNECTED_392, SV2V_UNCONNECTED_393, SV2V_UNCONNECTED_394, SV2V_UNCONNECTED_395, SV2V_UNCONNECTED_396, SV2V_UNCONNECTED_397, SV2V_UNCONNECTED_398, SV2V_UNCONNECTED_399, SV2V_UNCONNECTED_400, SV2V_UNCONNECTED_401, SV2V_UNCONNECTED_402, SV2V_UNCONNECTED_403, SV2V_UNCONNECTED_404, SV2V_UNCONNECTED_405, SV2V_UNCONNECTED_406, SV2V_UNCONNECTED_407, SV2V_UNCONNECTED_408, SV2V_UNCONNECTED_409, SV2V_UNCONNECTED_410, SV2V_UNCONNECTED_411, SV2V_UNCONNECTED_412, SV2V_UNCONNECTED_413, SV2V_UNCONNECTED_414, SV2V_UNCONNECTED_415, SV2V_UNCONNECTED_416, SV2V_UNCONNECTED_417, SV2V_UNCONNECTED_418, SV2V_UNCONNECTED_419, SV2V_UNCONNECTED_420, SV2V_UNCONNECTED_421, SV2V_UNCONNECTED_422, SV2V_UNCONNECTED_423, SV2V_UNCONNECTED_424, SV2V_UNCONNECTED_425, SV2V_UNCONNECTED_426, SV2V_UNCONNECTED_427, SV2V_UNCONNECTED_428, SV2V_UNCONNECTED_429, SV2V_UNCONNECTED_430, SV2V_UNCONNECTED_431, SV2V_UNCONNECTED_432, SV2V_UNCONNECTED_433, SV2V_UNCONNECTED_434, SV2V_UNCONNECTED_435, SV2V_UNCONNECTED_436, SV2V_UNCONNECTED_437, SV2V_UNCONNECTED_438, SV2V_UNCONNECTED_439, SV2V_UNCONNECTED_440, SV2V_UNCONNECTED_441, SV2V_UNCONNECTED_442, SV2V_UNCONNECTED_443, SV2V_UNCONNECTED_444, SV2V_UNCONNECTED_445, SV2V_UNCONNECTED_446, SV2V_UNCONNECTED_447, SV2V_UNCONNECTED_448, SV2V_UNCONNECTED_449, SV2V_UNCONNECTED_450, SV2V_UNCONNECTED_451, SV2V_UNCONNECTED_452, SV2V_UNCONNECTED_453, SV2V_UNCONNECTED_454, SV2V_UNCONNECTED_455, SV2V_UNCONNECTED_456, SV2V_UNCONNECTED_457, SV2V_UNCONNECTED_458, SV2V_UNCONNECTED_459, SV2V_UNCONNECTED_460, SV2V_UNCONNECTED_461, SV2V_UNCONNECTED_462, SV2V_UNCONNECTED_463, SV2V_UNCONNECTED_464, SV2V_UNCONNECTED_465, SV2V_UNCONNECTED_466, SV2V_UNCONNECTED_467, SV2V_UNCONNECTED_468, SV2V_UNCONNECTED_469, SV2V_UNCONNECTED_470, SV2V_UNCONNECTED_471, SV2V_UNCONNECTED_472, SV2V_UNCONNECTED_473, SV2V_UNCONNECTED_474, SV2V_UNCONNECTED_475, SV2V_UNCONNECTED_476, SV2V_UNCONNECTED_477, SV2V_UNCONNECTED_478, SV2V_UNCONNECTED_479, SV2V_UNCONNECTED_480, SV2V_UNCONNECTED_481, SV2V_UNCONNECTED_482, SV2V_UNCONNECTED_483, SV2V_UNCONNECTED_484, SV2V_UNCONNECTED_485, SV2V_UNCONNECTED_486, SV2V_UNCONNECTED_487, SV2V_UNCONNECTED_488, SV2V_UNCONNECTED_489, SV2V_UNCONNECTED_490, SV2V_UNCONNECTED_491, SV2V_UNCONNECTED_492, SV2V_UNCONNECTED_493, SV2V_UNCONNECTED_494, SV2V_UNCONNECTED_495, SV2V_UNCONNECTED_496, SV2V_UNCONNECTED_497, SV2V_UNCONNECTED_498, SV2V_UNCONNECTED_499, SV2V_UNCONNECTED_500, SV2V_UNCONNECTED_501, SV2V_UNCONNECTED_502, SV2V_UNCONNECTED_503, SV2V_UNCONNECTED_504, SV2V_UNCONNECTED_505, SV2V_UNCONNECTED_506, SV2V_UNCONNECTED_507, SV2V_UNCONNECTED_508, SV2V_UNCONNECTED_509, SV2V_UNCONNECTED_510, SV2V_UNCONNECTED_511, SV2V_UNCONNECTED_512, SV2V_UNCONNECTED_513, SV2V_UNCONNECTED_514, SV2V_UNCONNECTED_515, SV2V_UNCONNECTED_516, SV2V_UNCONNECTED_517, SV2V_UNCONNECTED_518, SV2V_UNCONNECTED_519, SV2V_UNCONNECTED_520, SV2V_UNCONNECTED_521, SV2V_UNCONNECTED_522, SV2V_UNCONNECTED_523, SV2V_UNCONNECTED_524, SV2V_UNCONNECTED_525, SV2V_UNCONNECTED_526, SV2V_UNCONNECTED_527, SV2V_UNCONNECTED_528, SV2V_UNCONNECTED_529, SV2V_UNCONNECTED_530, SV2V_UNCONNECTED_531, SV2V_UNCONNECTED_532, SV2V_UNCONNECTED_533, SV2V_UNCONNECTED_534, SV2V_UNCONNECTED_535, SV2V_UNCONNECTED_536, SV2V_UNCONNECTED_537, SV2V_UNCONNECTED_538, SV2V_UNCONNECTED_539, SV2V_UNCONNECTED_540, SV2V_UNCONNECTED_541, SV2V_UNCONNECTED_542, SV2V_UNCONNECTED_543, SV2V_UNCONNECTED_544, SV2V_UNCONNECTED_545, SV2V_UNCONNECTED_546, SV2V_UNCONNECTED_547, SV2V_UNCONNECTED_548, SV2V_UNCONNECTED_549, SV2V_UNCONNECTED_550, SV2V_UNCONNECTED_551, SV2V_UNCONNECTED_552, SV2V_UNCONNECTED_553, SV2V_UNCONNECTED_554, SV2V_UNCONNECTED_555, SV2V_UNCONNECTED_556, SV2V_UNCONNECTED_557, SV2V_UNCONNECTED_558, SV2V_UNCONNECTED_559, SV2V_UNCONNECTED_560, SV2V_UNCONNECTED_561, SV2V_UNCONNECTED_562, SV2V_UNCONNECTED_563, SV2V_UNCONNECTED_564, SV2V_UNCONNECTED_565, SV2V_UNCONNECTED_566, SV2V_UNCONNECTED_567, SV2V_UNCONNECTED_568, SV2V_UNCONNECTED_569, SV2V_UNCONNECTED_570, SV2V_UNCONNECTED_571, SV2V_UNCONNECTED_572, SV2V_UNCONNECTED_573, SV2V_UNCONNECTED_574, SV2V_UNCONNECTED_575, SV2V_UNCONNECTED_576, SV2V_UNCONNECTED_577, SV2V_UNCONNECTED_578, SV2V_UNCONNECTED_579, SV2V_UNCONNECTED_580, SV2V_UNCONNECTED_581, SV2V_UNCONNECTED_582, SV2V_UNCONNECTED_583, SV2V_UNCONNECTED_584, SV2V_UNCONNECTED_585, SV2V_UNCONNECTED_586, SV2V_UNCONNECTED_587, SV2V_UNCONNECTED_588, SV2V_UNCONNECTED_589, SV2V_UNCONNECTED_590, SV2V_UNCONNECTED_591, SV2V_UNCONNECTED_592, SV2V_UNCONNECTED_593, SV2V_UNCONNECTED_594, SV2V_UNCONNECTED_595, SV2V_UNCONNECTED_596, SV2V_UNCONNECTED_597, SV2V_UNCONNECTED_598, SV2V_UNCONNECTED_599, SV2V_UNCONNECTED_600, SV2V_UNCONNECTED_601, SV2V_UNCONNECTED_602, SV2V_UNCONNECTED_603, SV2V_UNCONNECTED_604, SV2V_UNCONNECTED_605, SV2V_UNCONNECTED_606, SV2V_UNCONNECTED_607, SV2V_UNCONNECTED_608, SV2V_UNCONNECTED_609, SV2V_UNCONNECTED_610, SV2V_UNCONNECTED_611, SV2V_UNCONNECTED_612, SV2V_UNCONNECTED_613, SV2V_UNCONNECTED_614, SV2V_UNCONNECTED_615, SV2V_UNCONNECTED_616, SV2V_UNCONNECTED_617, SV2V_UNCONNECTED_618, SV2V_UNCONNECTED_619, SV2V_UNCONNECTED_620, SV2V_UNCONNECTED_621, SV2V_UNCONNECTED_622, SV2V_UNCONNECTED_623, SV2V_UNCONNECTED_624, SV2V_UNCONNECTED_625, SV2V_UNCONNECTED_626, SV2V_UNCONNECTED_627, SV2V_UNCONNECTED_628, SV2V_UNCONNECTED_629, SV2V_UNCONNECTED_630, SV2V_UNCONNECTED_631, SV2V_UNCONNECTED_632, SV2V_UNCONNECTED_633, SV2V_UNCONNECTED_634, SV2V_UNCONNECTED_635, SV2V_UNCONNECTED_636, SV2V_UNCONNECTED_637, SV2V_UNCONNECTED_638, SV2V_UNCONNECTED_639, SV2V_UNCONNECTED_640, SV2V_UNCONNECTED_641, SV2V_UNCONNECTED_642, SV2V_UNCONNECTED_643, SV2V_UNCONNECTED_644, SV2V_UNCONNECTED_645, SV2V_UNCONNECTED_646, SV2V_UNCONNECTED_647, SV2V_UNCONNECTED_648, SV2V_UNCONNECTED_649, SV2V_UNCONNECTED_650, SV2V_UNCONNECTED_651, SV2V_UNCONNECTED_652, SV2V_UNCONNECTED_653, SV2V_UNCONNECTED_654, SV2V_UNCONNECTED_655, SV2V_UNCONNECTED_656, SV2V_UNCONNECTED_657, SV2V_UNCONNECTED_658, SV2V_UNCONNECTED_659, SV2V_UNCONNECTED_660, SV2V_UNCONNECTED_661, SV2V_UNCONNECTED_662, SV2V_UNCONNECTED_663, SV2V_UNCONNECTED_664, SV2V_UNCONNECTED_665, SV2V_UNCONNECTED_666, SV2V_UNCONNECTED_667, SV2V_UNCONNECTED_668, SV2V_UNCONNECTED_669, SV2V_UNCONNECTED_670, SV2V_UNCONNECTED_671, SV2V_UNCONNECTED_672, SV2V_UNCONNECTED_673, SV2V_UNCONNECTED_674, SV2V_UNCONNECTED_675, SV2V_UNCONNECTED_676, SV2V_UNCONNECTED_677, SV2V_UNCONNECTED_678, SV2V_UNCONNECTED_679, SV2V_UNCONNECTED_680, SV2V_UNCONNECTED_681, SV2V_UNCONNECTED_682, SV2V_UNCONNECTED_683, SV2V_UNCONNECTED_684, SV2V_UNCONNECTED_685, SV2V_UNCONNECTED_686, SV2V_UNCONNECTED_687, SV2V_UNCONNECTED_688, SV2V_UNCONNECTED_689, SV2V_UNCONNECTED_690, SV2V_UNCONNECTED_691, SV2V_UNCONNECTED_692, SV2V_UNCONNECTED_693, SV2V_UNCONNECTED_694, SV2V_UNCONNECTED_695, SV2V_UNCONNECTED_696, SV2V_UNCONNECTED_697, SV2V_UNCONNECTED_698, SV2V_UNCONNECTED_699, SV2V_UNCONNECTED_700, SV2V_UNCONNECTED_701, SV2V_UNCONNECTED_702, SV2V_UNCONNECTED_703, SV2V_UNCONNECTED_704, SV2V_UNCONNECTED_705, SV2V_UNCONNECTED_706, SV2V_UNCONNECTED_707, SV2V_UNCONNECTED_708, SV2V_UNCONNECTED_709, SV2V_UNCONNECTED_710, SV2V_UNCONNECTED_711, SV2V_UNCONNECTED_712, SV2V_UNCONNECTED_713, SV2V_UNCONNECTED_714, SV2V_UNCONNECTED_715, SV2V_UNCONNECTED_716, SV2V_UNCONNECTED_717, SV2V_UNCONNECTED_718, SV2V_UNCONNECTED_719, SV2V_UNCONNECTED_720, SV2V_UNCONNECTED_721, SV2V_UNCONNECTED_722, SV2V_UNCONNECTED_723, SV2V_UNCONNECTED_724, SV2V_UNCONNECTED_725, SV2V_UNCONNECTED_726, SV2V_UNCONNECTED_727, SV2V_UNCONNECTED_728, SV2V_UNCONNECTED_729, SV2V_UNCONNECTED_730, SV2V_UNCONNECTED_731, SV2V_UNCONNECTED_732, SV2V_UNCONNECTED_733, SV2V_UNCONNECTED_734, SV2V_UNCONNECTED_735, SV2V_UNCONNECTED_736, SV2V_UNCONNECTED_737, SV2V_UNCONNECTED_738, SV2V_UNCONNECTED_739, SV2V_UNCONNECTED_740, SV2V_UNCONNECTED_741, SV2V_UNCONNECTED_742, SV2V_UNCONNECTED_743, SV2V_UNCONNECTED_744, SV2V_UNCONNECTED_745, SV2V_UNCONNECTED_746, SV2V_UNCONNECTED_747, SV2V_UNCONNECTED_748, SV2V_UNCONNECTED_749, SV2V_UNCONNECTED_750, SV2V_UNCONNECTED_751, SV2V_UNCONNECTED_752, SV2V_UNCONNECTED_753, SV2V_UNCONNECTED_754, SV2V_UNCONNECTED_755, SV2V_UNCONNECTED_756, SV2V_UNCONNECTED_757, SV2V_UNCONNECTED_758, SV2V_UNCONNECTED_759, SV2V_UNCONNECTED_760, SV2V_UNCONNECTED_761, SV2V_UNCONNECTED_762, SV2V_UNCONNECTED_763, SV2V_UNCONNECTED_764, SV2V_UNCONNECTED_765, SV2V_UNCONNECTED_766, SV2V_UNCONNECTED_767, SV2V_UNCONNECTED_768, SV2V_UNCONNECTED_769, SV2V_UNCONNECTED_770, SV2V_UNCONNECTED_771, SV2V_UNCONNECTED_772, SV2V_UNCONNECTED_773, SV2V_UNCONNECTED_774, SV2V_UNCONNECTED_775, SV2V_UNCONNECTED_776, SV2V_UNCONNECTED_777, SV2V_UNCONNECTED_778, SV2V_UNCONNECTED_779, SV2V_UNCONNECTED_780, SV2V_UNCONNECTED_781, SV2V_UNCONNECTED_782, SV2V_UNCONNECTED_783, SV2V_UNCONNECTED_784, SV2V_UNCONNECTED_785, SV2V_UNCONNECTED_786, SV2V_UNCONNECTED_787, SV2V_UNCONNECTED_788, SV2V_UNCONNECTED_789, SV2V_UNCONNECTED_790, SV2V_UNCONNECTED_791, SV2V_UNCONNECTED_792, SV2V_UNCONNECTED_793, SV2V_UNCONNECTED_794, SV2V_UNCONNECTED_795, SV2V_UNCONNECTED_796, SV2V_UNCONNECTED_797, SV2V_UNCONNECTED_798, SV2V_UNCONNECTED_799, SV2V_UNCONNECTED_800, SV2V_UNCONNECTED_801, SV2V_UNCONNECTED_802, SV2V_UNCONNECTED_803, SV2V_UNCONNECTED_804, SV2V_UNCONNECTED_805, SV2V_UNCONNECTED_806, SV2V_UNCONNECTED_807, SV2V_UNCONNECTED_808, SV2V_UNCONNECTED_809, SV2V_UNCONNECTED_810, SV2V_UNCONNECTED_811, SV2V_UNCONNECTED_812, SV2V_UNCONNECTED_813, SV2V_UNCONNECTED_814, SV2V_UNCONNECTED_815, SV2V_UNCONNECTED_816, SV2V_UNCONNECTED_817, SV2V_UNCONNECTED_818, SV2V_UNCONNECTED_819, SV2V_UNCONNECTED_820, SV2V_UNCONNECTED_821, SV2V_UNCONNECTED_822, SV2V_UNCONNECTED_823, SV2V_UNCONNECTED_824, SV2V_UNCONNECTED_825, SV2V_UNCONNECTED_826, SV2V_UNCONNECTED_827, SV2V_UNCONNECTED_828, SV2V_UNCONNECTED_829, SV2V_UNCONNECTED_830, SV2V_UNCONNECTED_831, SV2V_UNCONNECTED_832, SV2V_UNCONNECTED_833, SV2V_UNCONNECTED_834, SV2V_UNCONNECTED_835, SV2V_UNCONNECTED_836, SV2V_UNCONNECTED_837, SV2V_UNCONNECTED_838, SV2V_UNCONNECTED_839, SV2V_UNCONNECTED_840, SV2V_UNCONNECTED_841, SV2V_UNCONNECTED_842, SV2V_UNCONNECTED_843, SV2V_UNCONNECTED_844, SV2V_UNCONNECTED_845, SV2V_UNCONNECTED_846, SV2V_UNCONNECTED_847, SV2V_UNCONNECTED_848, SV2V_UNCONNECTED_849, SV2V_UNCONNECTED_850, SV2V_UNCONNECTED_851, SV2V_UNCONNECTED_852, SV2V_UNCONNECTED_853, SV2V_UNCONNECTED_854, SV2V_UNCONNECTED_855, SV2V_UNCONNECTED_856, SV2V_UNCONNECTED_857, SV2V_UNCONNECTED_858, SV2V_UNCONNECTED_859, SV2V_UNCONNECTED_860, SV2V_UNCONNECTED_861, SV2V_UNCONNECTED_862, SV2V_UNCONNECTED_863, SV2V_UNCONNECTED_864, SV2V_UNCONNECTED_865, SV2V_UNCONNECTED_866, SV2V_UNCONNECTED_867, SV2V_UNCONNECTED_868, SV2V_UNCONNECTED_869, SV2V_UNCONNECTED_870, SV2V_UNCONNECTED_871, SV2V_UNCONNECTED_872, SV2V_UNCONNECTED_873, SV2V_UNCONNECTED_874, SV2V_UNCONNECTED_875, SV2V_UNCONNECTED_876, SV2V_UNCONNECTED_877, SV2V_UNCONNECTED_878, SV2V_UNCONNECTED_879, SV2V_UNCONNECTED_880, SV2V_UNCONNECTED_881, SV2V_UNCONNECTED_882, SV2V_UNCONNECTED_883, SV2V_UNCONNECTED_884, SV2V_UNCONNECTED_885, SV2V_UNCONNECTED_886, SV2V_UNCONNECTED_887, SV2V_UNCONNECTED_888, SV2V_UNCONNECTED_889, SV2V_UNCONNECTED_890, SV2V_UNCONNECTED_891, SV2V_UNCONNECTED_892, SV2V_UNCONNECTED_893, SV2V_UNCONNECTED_894, SV2V_UNCONNECTED_895, SV2V_UNCONNECTED_896, SV2V_UNCONNECTED_897, SV2V_UNCONNECTED_898, SV2V_UNCONNECTED_899, SV2V_UNCONNECTED_900, SV2V_UNCONNECTED_901, SV2V_UNCONNECTED_902, SV2V_UNCONNECTED_903, SV2V_UNCONNECTED_904, SV2V_UNCONNECTED_905, SV2V_UNCONNECTED_906, SV2V_UNCONNECTED_907, SV2V_UNCONNECTED_908, SV2V_UNCONNECTED_909, SV2V_UNCONNECTED_910, SV2V_UNCONNECTED_911, SV2V_UNCONNECTED_912, SV2V_UNCONNECTED_913, SV2V_UNCONNECTED_914, SV2V_UNCONNECTED_915, SV2V_UNCONNECTED_916, SV2V_UNCONNECTED_917, SV2V_UNCONNECTED_918, SV2V_UNCONNECTED_919, SV2V_UNCONNECTED_920, SV2V_UNCONNECTED_921, SV2V_UNCONNECTED_922, SV2V_UNCONNECTED_923, SV2V_UNCONNECTED_924, SV2V_UNCONNECTED_925, SV2V_UNCONNECTED_926, SV2V_UNCONNECTED_927, SV2V_UNCONNECTED_928, SV2V_UNCONNECTED_929, SV2V_UNCONNECTED_930, SV2V_UNCONNECTED_931, SV2V_UNCONNECTED_932, SV2V_UNCONNECTED_933, SV2V_UNCONNECTED_934, SV2V_UNCONNECTED_935, SV2V_UNCONNECTED_936, SV2V_UNCONNECTED_937, SV2V_UNCONNECTED_938, SV2V_UNCONNECTED_939, SV2V_UNCONNECTED_940, SV2V_UNCONNECTED_941, SV2V_UNCONNECTED_942, SV2V_UNCONNECTED_943, SV2V_UNCONNECTED_944, SV2V_UNCONNECTED_945, SV2V_UNCONNECTED_946, SV2V_UNCONNECTED_947, SV2V_UNCONNECTED_948, SV2V_UNCONNECTED_949, SV2V_UNCONNECTED_950, SV2V_UNCONNECTED_951, SV2V_UNCONNECTED_952, SV2V_UNCONNECTED_953, SV2V_UNCONNECTED_954, SV2V_UNCONNECTED_955, SV2V_UNCONNECTED_956, SV2V_UNCONNECTED_957, SV2V_UNCONNECTED_958, SV2V_UNCONNECTED_959, SV2V_UNCONNECTED_960, SV2V_UNCONNECTED_961, SV2V_UNCONNECTED_962, SV2V_UNCONNECTED_963, SV2V_UNCONNECTED_964, SV2V_UNCONNECTED_965, SV2V_UNCONNECTED_966, SV2V_UNCONNECTED_967, SV2V_UNCONNECTED_968, SV2V_UNCONNECTED_969, SV2V_UNCONNECTED_970, SV2V_UNCONNECTED_971, SV2V_UNCONNECTED_972, SV2V_UNCONNECTED_973, SV2V_UNCONNECTED_974, SV2V_UNCONNECTED_975, SV2V_UNCONNECTED_976, SV2V_UNCONNECTED_977, SV2V_UNCONNECTED_978, SV2V_UNCONNECTED_979, SV2V_UNCONNECTED_980, SV2V_UNCONNECTED_981, SV2V_UNCONNECTED_982, SV2V_UNCONNECTED_983, SV2V_UNCONNECTED_984, SV2V_UNCONNECTED_985, SV2V_UNCONNECTED_986, SV2V_UNCONNECTED_987, SV2V_UNCONNECTED_988, SV2V_UNCONNECTED_989, SV2V_UNCONNECTED_990, SV2V_UNCONNECTED_991, SV2V_UNCONNECTED_992, SV2V_UNCONNECTED_993, SV2V_UNCONNECTED_994, SV2V_UNCONNECTED_995, SV2V_UNCONNECTED_996, SV2V_UNCONNECTED_997, SV2V_UNCONNECTED_998, SV2V_UNCONNECTED_999, SV2V_UNCONNECTED_1000, SV2V_UNCONNECTED_1001, SV2V_UNCONNECTED_1002, SV2V_UNCONNECTED_1003, SV2V_UNCONNECTED_1004, SV2V_UNCONNECTED_1005, SV2V_UNCONNECTED_1006, SV2V_UNCONNECTED_1007, SV2V_UNCONNECTED_1008, SV2V_UNCONNECTED_1009, SV2V_UNCONNECTED_1010, SV2V_UNCONNECTED_1011, SV2V_UNCONNECTED_1012, SV2V_UNCONNECTED_1013, SV2V_UNCONNECTED_1014, SV2V_UNCONNECTED_1015, SV2V_UNCONNECTED_1016, SV2V_UNCONNECTED_1017, SV2V_UNCONNECTED_1018, SV2V_UNCONNECTED_1019, SV2V_UNCONNECTED_1020, SV2V_UNCONNECTED_1021, SV2V_UNCONNECTED_1022, SV2V_UNCONNECTED_1023, SV2V_UNCONNECTED_1024, SV2V_UNCONNECTED_1025, SV2V_UNCONNECTED_1026, SV2V_UNCONNECTED_1027, SV2V_UNCONNECTED_1028, SV2V_UNCONNECTED_1029, SV2V_UNCONNECTED_1030, SV2V_UNCONNECTED_1031, SV2V_UNCONNECTED_1032, SV2V_UNCONNECTED_1033, SV2V_UNCONNECTED_1034, SV2V_UNCONNECTED_1035, SV2V_UNCONNECTED_1036, SV2V_UNCONNECTED_1037, SV2V_UNCONNECTED_1038, SV2V_UNCONNECTED_1039, SV2V_UNCONNECTED_1040, SV2V_UNCONNECTED_1041, SV2V_UNCONNECTED_1042, SV2V_UNCONNECTED_1043, SV2V_UNCONNECTED_1044, SV2V_UNCONNECTED_1045, SV2V_UNCONNECTED_1046, SV2V_UNCONNECTED_1047, SV2V_UNCONNECTED_1048, SV2V_UNCONNECTED_1049, SV2V_UNCONNECTED_1050, SV2V_UNCONNECTED_1051, SV2V_UNCONNECTED_1052, SV2V_UNCONNECTED_1053, SV2V_UNCONNECTED_1054, SV2V_UNCONNECTED_1055, SV2V_UNCONNECTED_1056, SV2V_UNCONNECTED_1057, SV2V_UNCONNECTED_1058, SV2V_UNCONNECTED_1059, SV2V_UNCONNECTED_1060, SV2V_UNCONNECTED_1061, SV2V_UNCONNECTED_1062, SV2V_UNCONNECTED_1063, SV2V_UNCONNECTED_1064, SV2V_UNCONNECTED_1065, SV2V_UNCONNECTED_1066, SV2V_UNCONNECTED_1067, SV2V_UNCONNECTED_1068, SV2V_UNCONNECTED_1069, SV2V_UNCONNECTED_1070, SV2V_UNCONNECTED_1071, SV2V_UNCONNECTED_1072, SV2V_UNCONNECTED_1073, SV2V_UNCONNECTED_1074, SV2V_UNCONNECTED_1075, SV2V_UNCONNECTED_1076, SV2V_UNCONNECTED_1077, SV2V_UNCONNECTED_1078, SV2V_UNCONNECTED_1079, SV2V_UNCONNECTED_1080, SV2V_UNCONNECTED_1081, SV2V_UNCONNECTED_1082, SV2V_UNCONNECTED_1083, SV2V_UNCONNECTED_1084, SV2V_UNCONNECTED_1085, SV2V_UNCONNECTED_1086, SV2V_UNCONNECTED_1087, SV2V_UNCONNECTED_1088, SV2V_UNCONNECTED_1089, SV2V_UNCONNECTED_1090, SV2V_UNCONNECTED_1091, SV2V_UNCONNECTED_1092, SV2V_UNCONNECTED_1093, SV2V_UNCONNECTED_1094, SV2V_UNCONNECTED_1095, SV2V_UNCONNECTED_1096, SV2V_UNCONNECTED_1097, SV2V_UNCONNECTED_1098, SV2V_UNCONNECTED_1099, SV2V_UNCONNECTED_1100, SV2V_UNCONNECTED_1101, SV2V_UNCONNECTED_1102, SV2V_UNCONNECTED_1103, SV2V_UNCONNECTED_1104, SV2V_UNCONNECTED_1105, SV2V_UNCONNECTED_1106, SV2V_UNCONNECTED_1107, SV2V_UNCONNECTED_1108, SV2V_UNCONNECTED_1109, SV2V_UNCONNECTED_1110, SV2V_UNCONNECTED_1111, SV2V_UNCONNECTED_1112, SV2V_UNCONNECTED_1113, SV2V_UNCONNECTED_1114, SV2V_UNCONNECTED_1115, SV2V_UNCONNECTED_1116, SV2V_UNCONNECTED_1117, SV2V_UNCONNECTED_1118, SV2V_UNCONNECTED_1119, SV2V_UNCONNECTED_1120, SV2V_UNCONNECTED_1121, SV2V_UNCONNECTED_1122, SV2V_UNCONNECTED_1123, SV2V_UNCONNECTED_1124, SV2V_UNCONNECTED_1125, SV2V_UNCONNECTED_1126, SV2V_UNCONNECTED_1127, SV2V_UNCONNECTED_1128, SV2V_UNCONNECTED_1129, SV2V_UNCONNECTED_1130, SV2V_UNCONNECTED_1131, SV2V_UNCONNECTED_1132, SV2V_UNCONNECTED_1133, SV2V_UNCONNECTED_1134, SV2V_UNCONNECTED_1135, SV2V_UNCONNECTED_1136, SV2V_UNCONNECTED_1137, SV2V_UNCONNECTED_1138, SV2V_UNCONNECTED_1139, SV2V_UNCONNECTED_1140, SV2V_UNCONNECTED_1141, SV2V_UNCONNECTED_1142, SV2V_UNCONNECTED_1143, SV2V_UNCONNECTED_1144, SV2V_UNCONNECTED_1145, SV2V_UNCONNECTED_1146, SV2V_UNCONNECTED_1147, SV2V_UNCONNECTED_1148, SV2V_UNCONNECTED_1149, SV2V_UNCONNECTED_1150, SV2V_UNCONNECTED_1151, SV2V_UNCONNECTED_1152, SV2V_UNCONNECTED_1153, SV2V_UNCONNECTED_1154, SV2V_UNCONNECTED_1155, SV2V_UNCONNECTED_1156, SV2V_UNCONNECTED_1157, SV2V_UNCONNECTED_1158, SV2V_UNCONNECTED_1159, SV2V_UNCONNECTED_1160, SV2V_UNCONNECTED_1161, SV2V_UNCONNECTED_1162, SV2V_UNCONNECTED_1163, SV2V_UNCONNECTED_1164, SV2V_UNCONNECTED_1165, SV2V_UNCONNECTED_1166, SV2V_UNCONNECTED_1167, SV2V_UNCONNECTED_1168, SV2V_UNCONNECTED_1169, SV2V_UNCONNECTED_1170, SV2V_UNCONNECTED_1171, SV2V_UNCONNECTED_1172, SV2V_UNCONNECTED_1173, SV2V_UNCONNECTED_1174, SV2V_UNCONNECTED_1175, SV2V_UNCONNECTED_1176, SV2V_UNCONNECTED_1177, SV2V_UNCONNECTED_1178, SV2V_UNCONNECTED_1179, SV2V_UNCONNECTED_1180, SV2V_UNCONNECTED_1181, SV2V_UNCONNECTED_1182, SV2V_UNCONNECTED_1183, SV2V_UNCONNECTED_1184, SV2V_UNCONNECTED_1185, SV2V_UNCONNECTED_1186, SV2V_UNCONNECTED_1187, SV2V_UNCONNECTED_1188, SV2V_UNCONNECTED_1189, SV2V_UNCONNECTED_1190, SV2V_UNCONNECTED_1191, SV2V_UNCONNECTED_1192, SV2V_UNCONNECTED_1193, SV2V_UNCONNECTED_1194, SV2V_UNCONNECTED_1195, SV2V_UNCONNECTED_1196, SV2V_UNCONNECTED_1197, SV2V_UNCONNECTED_1198, SV2V_UNCONNECTED_1199, SV2V_UNCONNECTED_1200, SV2V_UNCONNECTED_1201, SV2V_UNCONNECTED_1202, SV2V_UNCONNECTED_1203, SV2V_UNCONNECTED_1204, SV2V_UNCONNECTED_1205, SV2V_UNCONNECTED_1206, SV2V_UNCONNECTED_1207, SV2V_UNCONNECTED_1208, SV2V_UNCONNECTED_1209, SV2V_UNCONNECTED_1210, SV2V_UNCONNECTED_1211, SV2V_UNCONNECTED_1212, SV2V_UNCONNECTED_1213, SV2V_UNCONNECTED_1214, SV2V_UNCONNECTED_1215, SV2V_UNCONNECTED_1216, SV2V_UNCONNECTED_1217, SV2V_UNCONNECTED_1218, SV2V_UNCONNECTED_1219, SV2V_UNCONNECTED_1220, SV2V_UNCONNECTED_1221, SV2V_UNCONNECTED_1222, SV2V_UNCONNECTED_1223, SV2V_UNCONNECTED_1224, SV2V_UNCONNECTED_1225, SV2V_UNCONNECTED_1226, SV2V_UNCONNECTED_1227, SV2V_UNCONNECTED_1228, SV2V_UNCONNECTED_1229, SV2V_UNCONNECTED_1230, SV2V_UNCONNECTED_1231, SV2V_UNCONNECTED_1232, SV2V_UNCONNECTED_1233, SV2V_UNCONNECTED_1234, SV2V_UNCONNECTED_1235, SV2V_UNCONNECTED_1236, SV2V_UNCONNECTED_1237, SV2V_UNCONNECTED_1238, SV2V_UNCONNECTED_1239, SV2V_UNCONNECTED_1240, SV2V_UNCONNECTED_1241, SV2V_UNCONNECTED_1242, SV2V_UNCONNECTED_1243, SV2V_UNCONNECTED_1244, SV2V_UNCONNECTED_1245, SV2V_UNCONNECTED_1246, SV2V_UNCONNECTED_1247, SV2V_UNCONNECTED_1248, SV2V_UNCONNECTED_1249, SV2V_UNCONNECTED_1250, SV2V_UNCONNECTED_1251, SV2V_UNCONNECTED_1252, SV2V_UNCONNECTED_1253, SV2V_UNCONNECTED_1254, SV2V_UNCONNECTED_1255, SV2V_UNCONNECTED_1256, SV2V_UNCONNECTED_1257, SV2V_UNCONNECTED_1258, SV2V_UNCONNECTED_1259, SV2V_UNCONNECTED_1260, SV2V_UNCONNECTED_1261, SV2V_UNCONNECTED_1262, SV2V_UNCONNECTED_1263, SV2V_UNCONNECTED_1264, SV2V_UNCONNECTED_1265, SV2V_UNCONNECTED_1266, SV2V_UNCONNECTED_1267, SV2V_UNCONNECTED_1268, SV2V_UNCONNECTED_1269, SV2V_UNCONNECTED_1270, SV2V_UNCONNECTED_1271, SV2V_UNCONNECTED_1272, SV2V_UNCONNECTED_1273, SV2V_UNCONNECTED_1274, SV2V_UNCONNECTED_1275, SV2V_UNCONNECTED_1276, SV2V_UNCONNECTED_1277, SV2V_UNCONNECTED_1278, SV2V_UNCONNECTED_1279, SV2V_UNCONNECTED_1280, SV2V_UNCONNECTED_1281, SV2V_UNCONNECTED_1282, SV2V_UNCONNECTED_1283, SV2V_UNCONNECTED_1284, SV2V_UNCONNECTED_1285, SV2V_UNCONNECTED_1286, SV2V_UNCONNECTED_1287, SV2V_UNCONNECTED_1288, SV2V_UNCONNECTED_1289, SV2V_UNCONNECTED_1290, SV2V_UNCONNECTED_1291, SV2V_UNCONNECTED_1292, SV2V_UNCONNECTED_1293, SV2V_UNCONNECTED_1294, SV2V_UNCONNECTED_1295, SV2V_UNCONNECTED_1296, SV2V_UNCONNECTED_1297, SV2V_UNCONNECTED_1298, SV2V_UNCONNECTED_1299, SV2V_UNCONNECTED_1300, SV2V_UNCONNECTED_1301, SV2V_UNCONNECTED_1302, SV2V_UNCONNECTED_1303, SV2V_UNCONNECTED_1304, SV2V_UNCONNECTED_1305, SV2V_UNCONNECTED_1306, SV2V_UNCONNECTED_1307, SV2V_UNCONNECTED_1308, SV2V_UNCONNECTED_1309, SV2V_UNCONNECTED_1310, SV2V_UNCONNECTED_1311, SV2V_UNCONNECTED_1312, SV2V_UNCONNECTED_1313, SV2V_UNCONNECTED_1314, SV2V_UNCONNECTED_1315, SV2V_UNCONNECTED_1316, SV2V_UNCONNECTED_1317, SV2V_UNCONNECTED_1318, SV2V_UNCONNECTED_1319, SV2V_UNCONNECTED_1320, SV2V_UNCONNECTED_1321, SV2V_UNCONNECTED_1322, SV2V_UNCONNECTED_1323, SV2V_UNCONNECTED_1324, SV2V_UNCONNECTED_1325, SV2V_UNCONNECTED_1326, SV2V_UNCONNECTED_1327, SV2V_UNCONNECTED_1328, SV2V_UNCONNECTED_1329, SV2V_UNCONNECTED_1330, SV2V_UNCONNECTED_1331, SV2V_UNCONNECTED_1332, SV2V_UNCONNECTED_1333, SV2V_UNCONNECTED_1334, SV2V_UNCONNECTED_1335, SV2V_UNCONNECTED_1336, SV2V_UNCONNECTED_1337, SV2V_UNCONNECTED_1338, SV2V_UNCONNECTED_1339, SV2V_UNCONNECTED_1340, SV2V_UNCONNECTED_1341, SV2V_UNCONNECTED_1342, SV2V_UNCONNECTED_1343, SV2V_UNCONNECTED_1344, SV2V_UNCONNECTED_1345, SV2V_UNCONNECTED_1346, SV2V_UNCONNECTED_1347, SV2V_UNCONNECTED_1348, SV2V_UNCONNECTED_1349, SV2V_UNCONNECTED_1350, SV2V_UNCONNECTED_1351, SV2V_UNCONNECTED_1352, SV2V_UNCONNECTED_1353, SV2V_UNCONNECTED_1354, SV2V_UNCONNECTED_1355, SV2V_UNCONNECTED_1356, SV2V_UNCONNECTED_1357, SV2V_UNCONNECTED_1358, SV2V_UNCONNECTED_1359, SV2V_UNCONNECTED_1360, SV2V_UNCONNECTED_1361, SV2V_UNCONNECTED_1362, SV2V_UNCONNECTED_1363, SV2V_UNCONNECTED_1364, SV2V_UNCONNECTED_1365, SV2V_UNCONNECTED_1366, SV2V_UNCONNECTED_1367, SV2V_UNCONNECTED_1368, SV2V_UNCONNECTED_1369, SV2V_UNCONNECTED_1370, SV2V_UNCONNECTED_1371, SV2V_UNCONNECTED_1372, SV2V_UNCONNECTED_1373, SV2V_UNCONNECTED_1374, SV2V_UNCONNECTED_1375, SV2V_UNCONNECTED_1376, SV2V_UNCONNECTED_1377, SV2V_UNCONNECTED_1378, SV2V_UNCONNECTED_1379, SV2V_UNCONNECTED_1380, SV2V_UNCONNECTED_1381, SV2V_UNCONNECTED_1382, SV2V_UNCONNECTED_1383, SV2V_UNCONNECTED_1384, SV2V_UNCONNECTED_1385, SV2V_UNCONNECTED_1386, SV2V_UNCONNECTED_1387, SV2V_UNCONNECTED_1388, SV2V_UNCONNECTED_1389, SV2V_UNCONNECTED_1390, SV2V_UNCONNECTED_1391, SV2V_UNCONNECTED_1392, SV2V_UNCONNECTED_1393, SV2V_UNCONNECTED_1394, SV2V_UNCONNECTED_1395, SV2V_UNCONNECTED_1396, SV2V_UNCONNECTED_1397, SV2V_UNCONNECTED_1398, SV2V_UNCONNECTED_1399, SV2V_UNCONNECTED_1400, SV2V_UNCONNECTED_1401, SV2V_UNCONNECTED_1402, SV2V_UNCONNECTED_1403, SV2V_UNCONNECTED_1404, SV2V_UNCONNECTED_1405, SV2V_UNCONNECTED_1406, SV2V_UNCONNECTED_1407, SV2V_UNCONNECTED_1408, SV2V_UNCONNECTED_1409, SV2V_UNCONNECTED_1410, SV2V_UNCONNECTED_1411, SV2V_UNCONNECTED_1412, SV2V_UNCONNECTED_1413, SV2V_UNCONNECTED_1414, SV2V_UNCONNECTED_1415, SV2V_UNCONNECTED_1416, SV2V_UNCONNECTED_1417, SV2V_UNCONNECTED_1418, SV2V_UNCONNECTED_1419, SV2V_UNCONNECTED_1420, SV2V_UNCONNECTED_1421, SV2V_UNCONNECTED_1422, SV2V_UNCONNECTED_1423, SV2V_UNCONNECTED_1424, SV2V_UNCONNECTED_1425, SV2V_UNCONNECTED_1426, SV2V_UNCONNECTED_1427, SV2V_UNCONNECTED_1428, SV2V_UNCONNECTED_1429, SV2V_UNCONNECTED_1430, SV2V_UNCONNECTED_1431, SV2V_UNCONNECTED_1432, SV2V_UNCONNECTED_1433, SV2V_UNCONNECTED_1434, SV2V_UNCONNECTED_1435, SV2V_UNCONNECTED_1436, SV2V_UNCONNECTED_1437, SV2V_UNCONNECTED_1438, SV2V_UNCONNECTED_1439, SV2V_UNCONNECTED_1440, SV2V_UNCONNECTED_1441, SV2V_UNCONNECTED_1442, SV2V_UNCONNECTED_1443, SV2V_UNCONNECTED_1444, SV2V_UNCONNECTED_1445, SV2V_UNCONNECTED_1446, SV2V_UNCONNECTED_1447, SV2V_UNCONNECTED_1448, SV2V_UNCONNECTED_1449, SV2V_UNCONNECTED_1450, SV2V_UNCONNECTED_1451, SV2V_UNCONNECTED_1452, SV2V_UNCONNECTED_1453, SV2V_UNCONNECTED_1454, SV2V_UNCONNECTED_1455, SV2V_UNCONNECTED_1456, SV2V_UNCONNECTED_1457, SV2V_UNCONNECTED_1458, SV2V_UNCONNECTED_1459, SV2V_UNCONNECTED_1460, SV2V_UNCONNECTED_1461, SV2V_UNCONNECTED_1462, SV2V_UNCONNECTED_1463, SV2V_UNCONNECTED_1464, SV2V_UNCONNECTED_1465, SV2V_UNCONNECTED_1466, SV2V_UNCONNECTED_1467, SV2V_UNCONNECTED_1468, SV2V_UNCONNECTED_1469, SV2V_UNCONNECTED_1470, SV2V_UNCONNECTED_1471, SV2V_UNCONNECTED_1472, SV2V_UNCONNECTED_1473, SV2V_UNCONNECTED_1474, SV2V_UNCONNECTED_1475, SV2V_UNCONNECTED_1476, SV2V_UNCONNECTED_1477, SV2V_UNCONNECTED_1478, SV2V_UNCONNECTED_1479, SV2V_UNCONNECTED_1480, SV2V_UNCONNECTED_1481, SV2V_UNCONNECTED_1482, SV2V_UNCONNECTED_1483, SV2V_UNCONNECTED_1484, SV2V_UNCONNECTED_1485, SV2V_UNCONNECTED_1486, SV2V_UNCONNECTED_1487, SV2V_UNCONNECTED_1488, SV2V_UNCONNECTED_1489, SV2V_UNCONNECTED_1490, SV2V_UNCONNECTED_1491, SV2V_UNCONNECTED_1492, SV2V_UNCONNECTED_1493, SV2V_UNCONNECTED_1494, SV2V_UNCONNECTED_1495, SV2V_UNCONNECTED_1496, SV2V_UNCONNECTED_1497, SV2V_UNCONNECTED_1498, SV2V_UNCONNECTED_1499, SV2V_UNCONNECTED_1500, SV2V_UNCONNECTED_1501, SV2V_UNCONNECTED_1502, SV2V_UNCONNECTED_1503, SV2V_UNCONNECTED_1504, SV2V_UNCONNECTED_1505, SV2V_UNCONNECTED_1506, SV2V_UNCONNECTED_1507, SV2V_UNCONNECTED_1508, SV2V_UNCONNECTED_1509, SV2V_UNCONNECTED_1510, SV2V_UNCONNECTED_1511, SV2V_UNCONNECTED_1512, SV2V_UNCONNECTED_1513, SV2V_UNCONNECTED_1514, SV2V_UNCONNECTED_1515, SV2V_UNCONNECTED_1516, SV2V_UNCONNECTED_1517, SV2V_UNCONNECTED_1518, SV2V_UNCONNECTED_1519, SV2V_UNCONNECTED_1520, SV2V_UNCONNECTED_1521, SV2V_UNCONNECTED_1522, SV2V_UNCONNECTED_1523, SV2V_UNCONNECTED_1524, SV2V_UNCONNECTED_1525, SV2V_UNCONNECTED_1526, SV2V_UNCONNECTED_1527, SV2V_UNCONNECTED_1528, SV2V_UNCONNECTED_1529, SV2V_UNCONNECTED_1530, SV2V_UNCONNECTED_1531, SV2V_UNCONNECTED_1532, SV2V_UNCONNECTED_1533, SV2V_UNCONNECTED_1534, SV2V_UNCONNECTED_1535, SV2V_UNCONNECTED_1536, SV2V_UNCONNECTED_1537, SV2V_UNCONNECTED_1538, SV2V_UNCONNECTED_1539, SV2V_UNCONNECTED_1540, SV2V_UNCONNECTED_1541, SV2V_UNCONNECTED_1542, SV2V_UNCONNECTED_1543, SV2V_UNCONNECTED_1544, SV2V_UNCONNECTED_1545, SV2V_UNCONNECTED_1546, SV2V_UNCONNECTED_1547, SV2V_UNCONNECTED_1548, SV2V_UNCONNECTED_1549, SV2V_UNCONNECTED_1550, SV2V_UNCONNECTED_1551, SV2V_UNCONNECTED_1552, SV2V_UNCONNECTED_1553, SV2V_UNCONNECTED_1554, SV2V_UNCONNECTED_1555, SV2V_UNCONNECTED_1556, SV2V_UNCONNECTED_1557, SV2V_UNCONNECTED_1558, SV2V_UNCONNECTED_1559, SV2V_UNCONNECTED_1560, SV2V_UNCONNECTED_1561, SV2V_UNCONNECTED_1562, SV2V_UNCONNECTED_1563, SV2V_UNCONNECTED_1564, SV2V_UNCONNECTED_1565, SV2V_UNCONNECTED_1566, SV2V_UNCONNECTED_1567, SV2V_UNCONNECTED_1568, SV2V_UNCONNECTED_1569, SV2V_UNCONNECTED_1570, SV2V_UNCONNECTED_1571, SV2V_UNCONNECTED_1572, SV2V_UNCONNECTED_1573, SV2V_UNCONNECTED_1574, SV2V_UNCONNECTED_1575, SV2V_UNCONNECTED_1576, SV2V_UNCONNECTED_1577, SV2V_UNCONNECTED_1578, SV2V_UNCONNECTED_1579, SV2V_UNCONNECTED_1580, SV2V_UNCONNECTED_1581, SV2V_UNCONNECTED_1582, SV2V_UNCONNECTED_1583, SV2V_UNCONNECTED_1584, SV2V_UNCONNECTED_1585, SV2V_UNCONNECTED_1586, SV2V_UNCONNECTED_1587, SV2V_UNCONNECTED_1588, SV2V_UNCONNECTED_1589, SV2V_UNCONNECTED_1590, SV2V_UNCONNECTED_1591, SV2V_UNCONNECTED_1592, SV2V_UNCONNECTED_1593, SV2V_UNCONNECTED_1594, SV2V_UNCONNECTED_1595, SV2V_UNCONNECTED_1596, SV2V_UNCONNECTED_1597, SV2V_UNCONNECTED_1598, SV2V_UNCONNECTED_1599, SV2V_UNCONNECTED_1600, SV2V_UNCONNECTED_1601, SV2V_UNCONNECTED_1602, SV2V_UNCONNECTED_1603, SV2V_UNCONNECTED_1604, SV2V_UNCONNECTED_1605, SV2V_UNCONNECTED_1606, SV2V_UNCONNECTED_1607, SV2V_UNCONNECTED_1608, SV2V_UNCONNECTED_1609, SV2V_UNCONNECTED_1610, SV2V_UNCONNECTED_1611, SV2V_UNCONNECTED_1612, SV2V_UNCONNECTED_1613, SV2V_UNCONNECTED_1614, SV2V_UNCONNECTED_1615, SV2V_UNCONNECTED_1616, SV2V_UNCONNECTED_1617, SV2V_UNCONNECTED_1618, SV2V_UNCONNECTED_1619, SV2V_UNCONNECTED_1620, SV2V_UNCONNECTED_1621, SV2V_UNCONNECTED_1622, SV2V_UNCONNECTED_1623, SV2V_UNCONNECTED_1624, SV2V_UNCONNECTED_1625, SV2V_UNCONNECTED_1626, SV2V_UNCONNECTED_1627, SV2V_UNCONNECTED_1628, SV2V_UNCONNECTED_1629, SV2V_UNCONNECTED_1630, SV2V_UNCONNECTED_1631, SV2V_UNCONNECTED_1632, SV2V_UNCONNECTED_1633, SV2V_UNCONNECTED_1634, SV2V_UNCONNECTED_1635, SV2V_UNCONNECTED_1636, SV2V_UNCONNECTED_1637, SV2V_UNCONNECTED_1638, SV2V_UNCONNECTED_1639, SV2V_UNCONNECTED_1640, SV2V_UNCONNECTED_1641, SV2V_UNCONNECTED_1642, SV2V_UNCONNECTED_1643, SV2V_UNCONNECTED_1644, SV2V_UNCONNECTED_1645, SV2V_UNCONNECTED_1646, SV2V_UNCONNECTED_1647, SV2V_UNCONNECTED_1648, SV2V_UNCONNECTED_1649, SV2V_UNCONNECTED_1650, SV2V_UNCONNECTED_1651, SV2V_UNCONNECTED_1652, SV2V_UNCONNECTED_1653, SV2V_UNCONNECTED_1654, SV2V_UNCONNECTED_1655, SV2V_UNCONNECTED_1656, SV2V_UNCONNECTED_1657, SV2V_UNCONNECTED_1658, SV2V_UNCONNECTED_1659, SV2V_UNCONNECTED_1660, SV2V_UNCONNECTED_1661, SV2V_UNCONNECTED_1662, SV2V_UNCONNECTED_1663, SV2V_UNCONNECTED_1664, SV2V_UNCONNECTED_1665, SV2V_UNCONNECTED_1666, SV2V_UNCONNECTED_1667, SV2V_UNCONNECTED_1668, SV2V_UNCONNECTED_1669, SV2V_UNCONNECTED_1670, SV2V_UNCONNECTED_1671, SV2V_UNCONNECTED_1672, SV2V_UNCONNECTED_1673, SV2V_UNCONNECTED_1674, SV2V_UNCONNECTED_1675, SV2V_UNCONNECTED_1676, SV2V_UNCONNECTED_1677, SV2V_UNCONNECTED_1678, SV2V_UNCONNECTED_1679, SV2V_UNCONNECTED_1680, SV2V_UNCONNECTED_1681, SV2V_UNCONNECTED_1682, SV2V_UNCONNECTED_1683, SV2V_UNCONNECTED_1684, SV2V_UNCONNECTED_1685, SV2V_UNCONNECTED_1686, SV2V_UNCONNECTED_1687, SV2V_UNCONNECTED_1688, SV2V_UNCONNECTED_1689, SV2V_UNCONNECTED_1690, SV2V_UNCONNECTED_1691, SV2V_UNCONNECTED_1692, SV2V_UNCONNECTED_1693, SV2V_UNCONNECTED_1694, SV2V_UNCONNECTED_1695, SV2V_UNCONNECTED_1696, SV2V_UNCONNECTED_1697, SV2V_UNCONNECTED_1698, SV2V_UNCONNECTED_1699, SV2V_UNCONNECTED_1700, SV2V_UNCONNECTED_1701, SV2V_UNCONNECTED_1702, SV2V_UNCONNECTED_1703, SV2V_UNCONNECTED_1704, SV2V_UNCONNECTED_1705, SV2V_UNCONNECTED_1706, SV2V_UNCONNECTED_1707, SV2V_UNCONNECTED_1708, SV2V_UNCONNECTED_1709, SV2V_UNCONNECTED_1710, SV2V_UNCONNECTED_1711, SV2V_UNCONNECTED_1712, SV2V_UNCONNECTED_1713, SV2V_UNCONNECTED_1714, SV2V_UNCONNECTED_1715, SV2V_UNCONNECTED_1716, SV2V_UNCONNECTED_1717, SV2V_UNCONNECTED_1718, SV2V_UNCONNECTED_1719, SV2V_UNCONNECTED_1720, SV2V_UNCONNECTED_1721, SV2V_UNCONNECTED_1722, SV2V_UNCONNECTED_1723, SV2V_UNCONNECTED_1724, SV2V_UNCONNECTED_1725, SV2V_UNCONNECTED_1726, SV2V_UNCONNECTED_1727, SV2V_UNCONNECTED_1728, SV2V_UNCONNECTED_1729, SV2V_UNCONNECTED_1730, SV2V_UNCONNECTED_1731, SV2V_UNCONNECTED_1732, SV2V_UNCONNECTED_1733, SV2V_UNCONNECTED_1734, SV2V_UNCONNECTED_1735, SV2V_UNCONNECTED_1736, SV2V_UNCONNECTED_1737, SV2V_UNCONNECTED_1738, SV2V_UNCONNECTED_1739, SV2V_UNCONNECTED_1740, SV2V_UNCONNECTED_1741, SV2V_UNCONNECTED_1742, SV2V_UNCONNECTED_1743, SV2V_UNCONNECTED_1744, SV2V_UNCONNECTED_1745, SV2V_UNCONNECTED_1746, SV2V_UNCONNECTED_1747, SV2V_UNCONNECTED_1748, SV2V_UNCONNECTED_1749, SV2V_UNCONNECTED_1750, SV2V_UNCONNECTED_1751, SV2V_UNCONNECTED_1752, SV2V_UNCONNECTED_1753, SV2V_UNCONNECTED_1754, SV2V_UNCONNECTED_1755, SV2V_UNCONNECTED_1756, SV2V_UNCONNECTED_1757, SV2V_UNCONNECTED_1758, SV2V_UNCONNECTED_1759, SV2V_UNCONNECTED_1760, SV2V_UNCONNECTED_1761, SV2V_UNCONNECTED_1762, SV2V_UNCONNECTED_1763, SV2V_UNCONNECTED_1764, SV2V_UNCONNECTED_1765, SV2V_UNCONNECTED_1766, SV2V_UNCONNECTED_1767, SV2V_UNCONNECTED_1768, SV2V_UNCONNECTED_1769, SV2V_UNCONNECTED_1770, SV2V_UNCONNECTED_1771, SV2V_UNCONNECTED_1772, SV2V_UNCONNECTED_1773, SV2V_UNCONNECTED_1774, SV2V_UNCONNECTED_1775, SV2V_UNCONNECTED_1776, SV2V_UNCONNECTED_1777, SV2V_UNCONNECTED_1778, SV2V_UNCONNECTED_1779, SV2V_UNCONNECTED_1780, SV2V_UNCONNECTED_1781, SV2V_UNCONNECTED_1782, SV2V_UNCONNECTED_1783, SV2V_UNCONNECTED_1784, SV2V_UNCONNECTED_1785, SV2V_UNCONNECTED_1786, SV2V_UNCONNECTED_1787, SV2V_UNCONNECTED_1788, SV2V_UNCONNECTED_1789, SV2V_UNCONNECTED_1790, SV2V_UNCONNECTED_1791, SV2V_UNCONNECTED_1792, SV2V_UNCONNECTED_1793, SV2V_UNCONNECTED_1794, SV2V_UNCONNECTED_1795, SV2V_UNCONNECTED_1796, SV2V_UNCONNECTED_1797, SV2V_UNCONNECTED_1798, SV2V_UNCONNECTED_1799, SV2V_UNCONNECTED_1800, SV2V_UNCONNECTED_1801, SV2V_UNCONNECTED_1802, SV2V_UNCONNECTED_1803, SV2V_UNCONNECTED_1804, SV2V_UNCONNECTED_1805, SV2V_UNCONNECTED_1806, SV2V_UNCONNECTED_1807, SV2V_UNCONNECTED_1808, SV2V_UNCONNECTED_1809, SV2V_UNCONNECTED_1810, SV2V_UNCONNECTED_1811, SV2V_UNCONNECTED_1812, SV2V_UNCONNECTED_1813, SV2V_UNCONNECTED_1814, SV2V_UNCONNECTED_1815, SV2V_UNCONNECTED_1816, SV2V_UNCONNECTED_1817, SV2V_UNCONNECTED_1818, SV2V_UNCONNECTED_1819, SV2V_UNCONNECTED_1820, SV2V_UNCONNECTED_1821, SV2V_UNCONNECTED_1822, SV2V_UNCONNECTED_1823, SV2V_UNCONNECTED_1824, SV2V_UNCONNECTED_1825, SV2V_UNCONNECTED_1826, SV2V_UNCONNECTED_1827, SV2V_UNCONNECTED_1828, SV2V_UNCONNECTED_1829, SV2V_UNCONNECTED_1830, SV2V_UNCONNECTED_1831, SV2V_UNCONNECTED_1832, SV2V_UNCONNECTED_1833, SV2V_UNCONNECTED_1834, SV2V_UNCONNECTED_1835, SV2V_UNCONNECTED_1836, SV2V_UNCONNECTED_1837, SV2V_UNCONNECTED_1838, SV2V_UNCONNECTED_1839, SV2V_UNCONNECTED_1840, SV2V_UNCONNECTED_1841, SV2V_UNCONNECTED_1842, SV2V_UNCONNECTED_1843, SV2V_UNCONNECTED_1844, SV2V_UNCONNECTED_1845, SV2V_UNCONNECTED_1846, SV2V_UNCONNECTED_1847, SV2V_UNCONNECTED_1848, SV2V_UNCONNECTED_1849, SV2V_UNCONNECTED_1850, SV2V_UNCONNECTED_1851, SV2V_UNCONNECTED_1852, SV2V_UNCONNECTED_1853, SV2V_UNCONNECTED_1854, SV2V_UNCONNECTED_1855, SV2V_UNCONNECTED_1856, SV2V_UNCONNECTED_1857, SV2V_UNCONNECTED_1858, SV2V_UNCONNECTED_1859, SV2V_UNCONNECTED_1860, SV2V_UNCONNECTED_1861, SV2V_UNCONNECTED_1862, SV2V_UNCONNECTED_1863, SV2V_UNCONNECTED_1864, SV2V_UNCONNECTED_1865, SV2V_UNCONNECTED_1866, SV2V_UNCONNECTED_1867, SV2V_UNCONNECTED_1868, SV2V_UNCONNECTED_1869, SV2V_UNCONNECTED_1870, SV2V_UNCONNECTED_1871, SV2V_UNCONNECTED_1872, SV2V_UNCONNECTED_1873, SV2V_UNCONNECTED_1874, SV2V_UNCONNECTED_1875, SV2V_UNCONNECTED_1876, SV2V_UNCONNECTED_1877, SV2V_UNCONNECTED_1878, SV2V_UNCONNECTED_1879, SV2V_UNCONNECTED_1880, SV2V_UNCONNECTED_1881, SV2V_UNCONNECTED_1882, SV2V_UNCONNECTED_1883, SV2V_UNCONNECTED_1884, SV2V_UNCONNECTED_1885, SV2V_UNCONNECTED_1886, SV2V_UNCONNECTED_1887, SV2V_UNCONNECTED_1888, SV2V_UNCONNECTED_1889, SV2V_UNCONNECTED_1890, SV2V_UNCONNECTED_1891, SV2V_UNCONNECTED_1892, SV2V_UNCONNECTED_1893, SV2V_UNCONNECTED_1894, SV2V_UNCONNECTED_1895, SV2V_UNCONNECTED_1896, SV2V_UNCONNECTED_1897, SV2V_UNCONNECTED_1898, SV2V_UNCONNECTED_1899, SV2V_UNCONNECTED_1900, SV2V_UNCONNECTED_1901, SV2V_UNCONNECTED_1902, SV2V_UNCONNECTED_1903, SV2V_UNCONNECTED_1904, SV2V_UNCONNECTED_1905, SV2V_UNCONNECTED_1906, SV2V_UNCONNECTED_1907, SV2V_UNCONNECTED_1908, SV2V_UNCONNECTED_1909, SV2V_UNCONNECTED_1910, SV2V_UNCONNECTED_1911, SV2V_UNCONNECTED_1912, SV2V_UNCONNECTED_1913, SV2V_UNCONNECTED_1914, SV2V_UNCONNECTED_1915, SV2V_UNCONNECTED_1916, SV2V_UNCONNECTED_1917, SV2V_UNCONNECTED_1918, SV2V_UNCONNECTED_1919, SV2V_UNCONNECTED_1920, SV2V_UNCONNECTED_1921, SV2V_UNCONNECTED_1922, SV2V_UNCONNECTED_1923, SV2V_UNCONNECTED_1924, SV2V_UNCONNECTED_1925, SV2V_UNCONNECTED_1926, SV2V_UNCONNECTED_1927, SV2V_UNCONNECTED_1928, SV2V_UNCONNECTED_1929, SV2V_UNCONNECTED_1930, SV2V_UNCONNECTED_1931, SV2V_UNCONNECTED_1932, SV2V_UNCONNECTED_1933, SV2V_UNCONNECTED_1934, SV2V_UNCONNECTED_1935, SV2V_UNCONNECTED_1936, SV2V_UNCONNECTED_1937, SV2V_UNCONNECTED_1938, SV2V_UNCONNECTED_1939, SV2V_UNCONNECTED_1940, SV2V_UNCONNECTED_1941, SV2V_UNCONNECTED_1942, SV2V_UNCONNECTED_1943, SV2V_UNCONNECTED_1944, SV2V_UNCONNECTED_1945, SV2V_UNCONNECTED_1946, SV2V_UNCONNECTED_1947, SV2V_UNCONNECTED_1948, SV2V_UNCONNECTED_1949, SV2V_UNCONNECTED_1950, SV2V_UNCONNECTED_1951, SV2V_UNCONNECTED_1952, SV2V_UNCONNECTED_1953, SV2V_UNCONNECTED_1954, SV2V_UNCONNECTED_1955, SV2V_UNCONNECTED_1956, SV2V_UNCONNECTED_1957, SV2V_UNCONNECTED_1958, SV2V_UNCONNECTED_1959, SV2V_UNCONNECTED_1960, SV2V_UNCONNECTED_1961, SV2V_UNCONNECTED_1962, SV2V_UNCONNECTED_1963, SV2V_UNCONNECTED_1964, SV2V_UNCONNECTED_1965, SV2V_UNCONNECTED_1966, SV2V_UNCONNECTED_1967, SV2V_UNCONNECTED_1968, SV2V_UNCONNECTED_1969, SV2V_UNCONNECTED_1970, SV2V_UNCONNECTED_1971, SV2V_UNCONNECTED_1972, SV2V_UNCONNECTED_1973, SV2V_UNCONNECTED_1974, SV2V_UNCONNECTED_1975, SV2V_UNCONNECTED_1976, SV2V_UNCONNECTED_1977, SV2V_UNCONNECTED_1978, SV2V_UNCONNECTED_1979, SV2V_UNCONNECTED_1980, SV2V_UNCONNECTED_1981, SV2V_UNCONNECTED_1982, SV2V_UNCONNECTED_1983, SV2V_UNCONNECTED_1984, SV2V_UNCONNECTED_1985, SV2V_UNCONNECTED_1986, SV2V_UNCONNECTED_1987, SV2V_UNCONNECTED_1988, SV2V_UNCONNECTED_1989, SV2V_UNCONNECTED_1990, SV2V_UNCONNECTED_1991, SV2V_UNCONNECTED_1992, SV2V_UNCONNECTED_1993, SV2V_UNCONNECTED_1994, SV2V_UNCONNECTED_1995, SV2V_UNCONNECTED_1996, SV2V_UNCONNECTED_1997, SV2V_UNCONNECTED_1998, SV2V_UNCONNECTED_1999, SV2V_UNCONNECTED_2000, SV2V_UNCONNECTED_2001, SV2V_UNCONNECTED_2002, SV2V_UNCONNECTED_2003, SV2V_UNCONNECTED_2004, SV2V_UNCONNECTED_2005, SV2V_UNCONNECTED_2006, SV2V_UNCONNECTED_2007, SV2V_UNCONNECTED_2008, SV2V_UNCONNECTED_2009, SV2V_UNCONNECTED_2010, SV2V_UNCONNECTED_2011, SV2V_UNCONNECTED_2012, SV2V_UNCONNECTED_2013, SV2V_UNCONNECTED_2014, SV2V_UNCONNECTED_2015, SV2V_UNCONNECTED_2016, SV2V_UNCONNECTED_2017, SV2V_UNCONNECTED_2018, SV2V_UNCONNECTED_2019, SV2V_UNCONNECTED_2020, SV2V_UNCONNECTED_2021, SV2V_UNCONNECTED_2022, SV2V_UNCONNECTED_2023, SV2V_UNCONNECTED_2024, SV2V_UNCONNECTED_2025, SV2V_UNCONNECTED_2026, SV2V_UNCONNECTED_2027, SV2V_UNCONNECTED_2028, SV2V_UNCONNECTED_2029, SV2V_UNCONNECTED_2030, SV2V_UNCONNECTED_2031, SV2V_UNCONNECTED_2032, SV2V_UNCONNECTED_2033, SV2V_UNCONNECTED_2034, SV2V_UNCONNECTED_2035, SV2V_UNCONNECTED_2036, SV2V_UNCONNECTED_2037, SV2V_UNCONNECTED_2038, SV2V_UNCONNECTED_2039, SV2V_UNCONNECTED_2040, SV2V_UNCONNECTED_2041, SV2V_UNCONNECTED_2042, SV2V_UNCONNECTED_2043, SV2V_UNCONNECTED_2044, SV2V_UNCONNECTED_2045, SV2V_UNCONNECTED_2046, SV2V_UNCONNECTED_2047, SV2V_UNCONNECTED_2048, SV2V_UNCONNECTED_2049, SV2V_UNCONNECTED_2050, SV2V_UNCONNECTED_2051, SV2V_UNCONNECTED_2052, SV2V_UNCONNECTED_2053, SV2V_UNCONNECTED_2054, SV2V_UNCONNECTED_2055, SV2V_UNCONNECTED_2056, SV2V_UNCONNECTED_2057, SV2V_UNCONNECTED_2058, SV2V_UNCONNECTED_2059, SV2V_UNCONNECTED_2060, SV2V_UNCONNECTED_2061, SV2V_UNCONNECTED_2062, SV2V_UNCONNECTED_2063, SV2V_UNCONNECTED_2064, SV2V_UNCONNECTED_2065, SV2V_UNCONNECTED_2066, SV2V_UNCONNECTED_2067, SV2V_UNCONNECTED_2068, SV2V_UNCONNECTED_2069, SV2V_UNCONNECTED_2070, SV2V_UNCONNECTED_2071, SV2V_UNCONNECTED_2072, SV2V_UNCONNECTED_2073, SV2V_UNCONNECTED_2074, SV2V_UNCONNECTED_2075, SV2V_UNCONNECTED_2076, SV2V_UNCONNECTED_2077, SV2V_UNCONNECTED_2078, SV2V_UNCONNECTED_2079, SV2V_UNCONNECTED_2080, SV2V_UNCONNECTED_2081, SV2V_UNCONNECTED_2082, SV2V_UNCONNECTED_2083, SV2V_UNCONNECTED_2084, SV2V_UNCONNECTED_2085, SV2V_UNCONNECTED_2086, SV2V_UNCONNECTED_2087, SV2V_UNCONNECTED_2088, SV2V_UNCONNECTED_2089, SV2V_UNCONNECTED_2090, SV2V_UNCONNECTED_2091, SV2V_UNCONNECTED_2092, SV2V_UNCONNECTED_2093, SV2V_UNCONNECTED_2094, SV2V_UNCONNECTED_2095, SV2V_UNCONNECTED_2096, SV2V_UNCONNECTED_2097, SV2V_UNCONNECTED_2098, SV2V_UNCONNECTED_2099, SV2V_UNCONNECTED_2100, SV2V_UNCONNECTED_2101, SV2V_UNCONNECTED_2102, SV2V_UNCONNECTED_2103, SV2V_UNCONNECTED_2104, SV2V_UNCONNECTED_2105, SV2V_UNCONNECTED_2106, SV2V_UNCONNECTED_2107, SV2V_UNCONNECTED_2108, SV2V_UNCONNECTED_2109, SV2V_UNCONNECTED_2110, SV2V_UNCONNECTED_2111, SV2V_UNCONNECTED_2112, SV2V_UNCONNECTED_2113, SV2V_UNCONNECTED_2114, SV2V_UNCONNECTED_2115, SV2V_UNCONNECTED_2116, SV2V_UNCONNECTED_2117, SV2V_UNCONNECTED_2118, SV2V_UNCONNECTED_2119, SV2V_UNCONNECTED_2120, SV2V_UNCONNECTED_2121, SV2V_UNCONNECTED_2122, SV2V_UNCONNECTED_2123, SV2V_UNCONNECTED_2124, SV2V_UNCONNECTED_2125, SV2V_UNCONNECTED_2126, SV2V_UNCONNECTED_2127, SV2V_UNCONNECTED_2128, SV2V_UNCONNECTED_2129, SV2V_UNCONNECTED_2130, SV2V_UNCONNECTED_2131, SV2V_UNCONNECTED_2132, SV2V_UNCONNECTED_2133, SV2V_UNCONNECTED_2134, SV2V_UNCONNECTED_2135, SV2V_UNCONNECTED_2136, SV2V_UNCONNECTED_2137, SV2V_UNCONNECTED_2138, SV2V_UNCONNECTED_2139, SV2V_UNCONNECTED_2140, SV2V_UNCONNECTED_2141, SV2V_UNCONNECTED_2142, SV2V_UNCONNECTED_2143, SV2V_UNCONNECTED_2144, SV2V_UNCONNECTED_2145, SV2V_UNCONNECTED_2146, SV2V_UNCONNECTED_2147, SV2V_UNCONNECTED_2148, SV2V_UNCONNECTED_2149, SV2V_UNCONNECTED_2150, SV2V_UNCONNECTED_2151, SV2V_UNCONNECTED_2152, SV2V_UNCONNECTED_2153, SV2V_UNCONNECTED_2154, SV2V_UNCONNECTED_2155, SV2V_UNCONNECTED_2156, SV2V_UNCONNECTED_2157, SV2V_UNCONNECTED_2158, SV2V_UNCONNECTED_2159, SV2V_UNCONNECTED_2160, SV2V_UNCONNECTED_2161, SV2V_UNCONNECTED_2162, SV2V_UNCONNECTED_2163, SV2V_UNCONNECTED_2164, SV2V_UNCONNECTED_2165, SV2V_UNCONNECTED_2166, SV2V_UNCONNECTED_2167, SV2V_UNCONNECTED_2168, SV2V_UNCONNECTED_2169, SV2V_UNCONNECTED_2170, SV2V_UNCONNECTED_2171, SV2V_UNCONNECTED_2172, SV2V_UNCONNECTED_2173, SV2V_UNCONNECTED_2174, SV2V_UNCONNECTED_2175, SV2V_UNCONNECTED_2176, SV2V_UNCONNECTED_2177, SV2V_UNCONNECTED_2178, SV2V_UNCONNECTED_2179, SV2V_UNCONNECTED_2180, SV2V_UNCONNECTED_2181, SV2V_UNCONNECTED_2182, SV2V_UNCONNECTED_2183, SV2V_UNCONNECTED_2184, SV2V_UNCONNECTED_2185, SV2V_UNCONNECTED_2186, SV2V_UNCONNECTED_2187, SV2V_UNCONNECTED_2188, SV2V_UNCONNECTED_2189, SV2V_UNCONNECTED_2190, SV2V_UNCONNECTED_2191, SV2V_UNCONNECTED_2192, SV2V_UNCONNECTED_2193, SV2V_UNCONNECTED_2194, SV2V_UNCONNECTED_2195, SV2V_UNCONNECTED_2196, SV2V_UNCONNECTED_2197, SV2V_UNCONNECTED_2198, SV2V_UNCONNECTED_2199, SV2V_UNCONNECTED_2200, SV2V_UNCONNECTED_2201, SV2V_UNCONNECTED_2202, SV2V_UNCONNECTED_2203, SV2V_UNCONNECTED_2204, SV2V_UNCONNECTED_2205, SV2V_UNCONNECTED_2206, SV2V_UNCONNECTED_2207, SV2V_UNCONNECTED_2208, SV2V_UNCONNECTED_2209, SV2V_UNCONNECTED_2210, SV2V_UNCONNECTED_2211, SV2V_UNCONNECTED_2212, SV2V_UNCONNECTED_2213, SV2V_UNCONNECTED_2214, SV2V_UNCONNECTED_2215, SV2V_UNCONNECTED_2216, SV2V_UNCONNECTED_2217, SV2V_UNCONNECTED_2218, SV2V_UNCONNECTED_2219, SV2V_UNCONNECTED_2220, SV2V_UNCONNECTED_2221, SV2V_UNCONNECTED_2222, SV2V_UNCONNECTED_2223, SV2V_UNCONNECTED_2224, SV2V_UNCONNECTED_2225, SV2V_UNCONNECTED_2226, SV2V_UNCONNECTED_2227, SV2V_UNCONNECTED_2228, SV2V_UNCONNECTED_2229, SV2V_UNCONNECTED_2230, SV2V_UNCONNECTED_2231, SV2V_UNCONNECTED_2232, SV2V_UNCONNECTED_2233, SV2V_UNCONNECTED_2234, SV2V_UNCONNECTED_2235, SV2V_UNCONNECTED_2236, SV2V_UNCONNECTED_2237, SV2V_UNCONNECTED_2238, SV2V_UNCONNECTED_2239, SV2V_UNCONNECTED_2240, SV2V_UNCONNECTED_2241, SV2V_UNCONNECTED_2242, SV2V_UNCONNECTED_2243, SV2V_UNCONNECTED_2244, SV2V_UNCONNECTED_2245, SV2V_UNCONNECTED_2246, SV2V_UNCONNECTED_2247, SV2V_UNCONNECTED_2248, SV2V_UNCONNECTED_2249, SV2V_UNCONNECTED_2250, SV2V_UNCONNECTED_2251, SV2V_UNCONNECTED_2252, SV2V_UNCONNECTED_2253, SV2V_UNCONNECTED_2254, SV2V_UNCONNECTED_2255, SV2V_UNCONNECTED_2256, SV2V_UNCONNECTED_2257, SV2V_UNCONNECTED_2258, SV2V_UNCONNECTED_2259, SV2V_UNCONNECTED_2260, SV2V_UNCONNECTED_2261, SV2V_UNCONNECTED_2262, SV2V_UNCONNECTED_2263, SV2V_UNCONNECTED_2264, SV2V_UNCONNECTED_2265, SV2V_UNCONNECTED_2266, SV2V_UNCONNECTED_2267, SV2V_UNCONNECTED_2268, SV2V_UNCONNECTED_2269, SV2V_UNCONNECTED_2270, SV2V_UNCONNECTED_2271, SV2V_UNCONNECTED_2272, SV2V_UNCONNECTED_2273, SV2V_UNCONNECTED_2274, SV2V_UNCONNECTED_2275, SV2V_UNCONNECTED_2276, SV2V_UNCONNECTED_2277, SV2V_UNCONNECTED_2278, SV2V_UNCONNECTED_2279, SV2V_UNCONNECTED_2280, SV2V_UNCONNECTED_2281, SV2V_UNCONNECTED_2282, SV2V_UNCONNECTED_2283, SV2V_UNCONNECTED_2284, SV2V_UNCONNECTED_2285, SV2V_UNCONNECTED_2286, SV2V_UNCONNECTED_2287, SV2V_UNCONNECTED_2288, SV2V_UNCONNECTED_2289, SV2V_UNCONNECTED_2290, SV2V_UNCONNECTED_2291, SV2V_UNCONNECTED_2292, SV2V_UNCONNECTED_2293, SV2V_UNCONNECTED_2294, SV2V_UNCONNECTED_2295, SV2V_UNCONNECTED_2296, SV2V_UNCONNECTED_2297, SV2V_UNCONNECTED_2298, SV2V_UNCONNECTED_2299, SV2V_UNCONNECTED_2300, SV2V_UNCONNECTED_2301, SV2V_UNCONNECTED_2302, SV2V_UNCONNECTED_2303, SV2V_UNCONNECTED_2304, SV2V_UNCONNECTED_2305, SV2V_UNCONNECTED_2306, SV2V_UNCONNECTED_2307, SV2V_UNCONNECTED_2308, SV2V_UNCONNECTED_2309, SV2V_UNCONNECTED_2310, SV2V_UNCONNECTED_2311, SV2V_UNCONNECTED_2312, SV2V_UNCONNECTED_2313, SV2V_UNCONNECTED_2314, SV2V_UNCONNECTED_2315, SV2V_UNCONNECTED_2316, SV2V_UNCONNECTED_2317, SV2V_UNCONNECTED_2318, SV2V_UNCONNECTED_2319, SV2V_UNCONNECTED_2320, SV2V_UNCONNECTED_2321, SV2V_UNCONNECTED_2322, SV2V_UNCONNECTED_2323, SV2V_UNCONNECTED_2324, SV2V_UNCONNECTED_2325, SV2V_UNCONNECTED_2326, SV2V_UNCONNECTED_2327, SV2V_UNCONNECTED_2328, SV2V_UNCONNECTED_2329, SV2V_UNCONNECTED_2330, SV2V_UNCONNECTED_2331, SV2V_UNCONNECTED_2332, SV2V_UNCONNECTED_2333, SV2V_UNCONNECTED_2334, SV2V_UNCONNECTED_2335, SV2V_UNCONNECTED_2336, SV2V_UNCONNECTED_2337, SV2V_UNCONNECTED_2338, SV2V_UNCONNECTED_2339, SV2V_UNCONNECTED_2340, SV2V_UNCONNECTED_2341, SV2V_UNCONNECTED_2342, SV2V_UNCONNECTED_2343, SV2V_UNCONNECTED_2344, SV2V_UNCONNECTED_2345, SV2V_UNCONNECTED_2346, SV2V_UNCONNECTED_2347, SV2V_UNCONNECTED_2348, SV2V_UNCONNECTED_2349, SV2V_UNCONNECTED_2350, SV2V_UNCONNECTED_2351, SV2V_UNCONNECTED_2352, SV2V_UNCONNECTED_2353, SV2V_UNCONNECTED_2354, SV2V_UNCONNECTED_2355, SV2V_UNCONNECTED_2356, SV2V_UNCONNECTED_2357, SV2V_UNCONNECTED_2358, SV2V_UNCONNECTED_2359, SV2V_UNCONNECTED_2360, SV2V_UNCONNECTED_2361, SV2V_UNCONNECTED_2362, SV2V_UNCONNECTED_2363, SV2V_UNCONNECTED_2364, SV2V_UNCONNECTED_2365, SV2V_UNCONNECTED_2366, SV2V_UNCONNECTED_2367, SV2V_UNCONNECTED_2368, SV2V_UNCONNECTED_2369, SV2V_UNCONNECTED_2370, SV2V_UNCONNECTED_2371, SV2V_UNCONNECTED_2372, SV2V_UNCONNECTED_2373, SV2V_UNCONNECTED_2374, SV2V_UNCONNECTED_2375, SV2V_UNCONNECTED_2376, SV2V_UNCONNECTED_2377, SV2V_UNCONNECTED_2378, SV2V_UNCONNECTED_2379, SV2V_UNCONNECTED_2380, SV2V_UNCONNECTED_2381, SV2V_UNCONNECTED_2382, SV2V_UNCONNECTED_2383, SV2V_UNCONNECTED_2384, SV2V_UNCONNECTED_2385, SV2V_UNCONNECTED_2386, SV2V_UNCONNECTED_2387, SV2V_UNCONNECTED_2388, SV2V_UNCONNECTED_2389, SV2V_UNCONNECTED_2390, SV2V_UNCONNECTED_2391, SV2V_UNCONNECTED_2392, SV2V_UNCONNECTED_2393, SV2V_UNCONNECTED_2394, SV2V_UNCONNECTED_2395, SV2V_UNCONNECTED_2396, SV2V_UNCONNECTED_2397, SV2V_UNCONNECTED_2398, SV2V_UNCONNECTED_2399, SV2V_UNCONNECTED_2400, SV2V_UNCONNECTED_2401, SV2V_UNCONNECTED_2402, SV2V_UNCONNECTED_2403, SV2V_UNCONNECTED_2404, SV2V_UNCONNECTED_2405, SV2V_UNCONNECTED_2406, SV2V_UNCONNECTED_2407, SV2V_UNCONNECTED_2408, SV2V_UNCONNECTED_2409, SV2V_UNCONNECTED_2410, SV2V_UNCONNECTED_2411, SV2V_UNCONNECTED_2412, SV2V_UNCONNECTED_2413, SV2V_UNCONNECTED_2414, SV2V_UNCONNECTED_2415, SV2V_UNCONNECTED_2416, SV2V_UNCONNECTED_2417, SV2V_UNCONNECTED_2418, SV2V_UNCONNECTED_2419, SV2V_UNCONNECTED_2420, SV2V_UNCONNECTED_2421, SV2V_UNCONNECTED_2422, SV2V_UNCONNECTED_2423, SV2V_UNCONNECTED_2424, SV2V_UNCONNECTED_2425, SV2V_UNCONNECTED_2426, SV2V_UNCONNECTED_2427, SV2V_UNCONNECTED_2428, SV2V_UNCONNECTED_2429, SV2V_UNCONNECTED_2430, SV2V_UNCONNECTED_2431, SV2V_UNCONNECTED_2432, SV2V_UNCONNECTED_2433, SV2V_UNCONNECTED_2434, SV2V_UNCONNECTED_2435, SV2V_UNCONNECTED_2436, SV2V_UNCONNECTED_2437, SV2V_UNCONNECTED_2438, SV2V_UNCONNECTED_2439, SV2V_UNCONNECTED_2440, SV2V_UNCONNECTED_2441, SV2V_UNCONNECTED_2442, SV2V_UNCONNECTED_2443, SV2V_UNCONNECTED_2444, SV2V_UNCONNECTED_2445, SV2V_UNCONNECTED_2446, SV2V_UNCONNECTED_2447, SV2V_UNCONNECTED_2448, SV2V_UNCONNECTED_2449, SV2V_UNCONNECTED_2450, SV2V_UNCONNECTED_2451, SV2V_UNCONNECTED_2452, SV2V_UNCONNECTED_2453, SV2V_UNCONNECTED_2454, SV2V_UNCONNECTED_2455, SV2V_UNCONNECTED_2456, SV2V_UNCONNECTED_2457, SV2V_UNCONNECTED_2458, SV2V_UNCONNECTED_2459, SV2V_UNCONNECTED_2460, SV2V_UNCONNECTED_2461, SV2V_UNCONNECTED_2462, SV2V_UNCONNECTED_2463, SV2V_UNCONNECTED_2464, SV2V_UNCONNECTED_2465, SV2V_UNCONNECTED_2466, SV2V_UNCONNECTED_2467, SV2V_UNCONNECTED_2468, SV2V_UNCONNECTED_2469, SV2V_UNCONNECTED_2470, SV2V_UNCONNECTED_2471, SV2V_UNCONNECTED_2472, SV2V_UNCONNECTED_2473, SV2V_UNCONNECTED_2474, SV2V_UNCONNECTED_2475, SV2V_UNCONNECTED_2476, SV2V_UNCONNECTED_2477, SV2V_UNCONNECTED_2478, SV2V_UNCONNECTED_2479, SV2V_UNCONNECTED_2480, SV2V_UNCONNECTED_2481, SV2V_UNCONNECTED_2482, SV2V_UNCONNECTED_2483, SV2V_UNCONNECTED_2484, SV2V_UNCONNECTED_2485, SV2V_UNCONNECTED_2486, SV2V_UNCONNECTED_2487, SV2V_UNCONNECTED_2488, SV2V_UNCONNECTED_2489, SV2V_UNCONNECTED_2490, SV2V_UNCONNECTED_2491, SV2V_UNCONNECTED_2492, SV2V_UNCONNECTED_2493, SV2V_UNCONNECTED_2494, SV2V_UNCONNECTED_2495, SV2V_UNCONNECTED_2496, SV2V_UNCONNECTED_2497, SV2V_UNCONNECTED_2498, SV2V_UNCONNECTED_2499, SV2V_UNCONNECTED_2500, SV2V_UNCONNECTED_2501, SV2V_UNCONNECTED_2502, SV2V_UNCONNECTED_2503, SV2V_UNCONNECTED_2504, SV2V_UNCONNECTED_2505, SV2V_UNCONNECTED_2506, SV2V_UNCONNECTED_2507, SV2V_UNCONNECTED_2508, SV2V_UNCONNECTED_2509, SV2V_UNCONNECTED_2510, SV2V_UNCONNECTED_2511, SV2V_UNCONNECTED_2512, SV2V_UNCONNECTED_2513, SV2V_UNCONNECTED_2514, SV2V_UNCONNECTED_2515, SV2V_UNCONNECTED_2516, SV2V_UNCONNECTED_2517, SV2V_UNCONNECTED_2518, SV2V_UNCONNECTED_2519, SV2V_UNCONNECTED_2520, SV2V_UNCONNECTED_2521, SV2V_UNCONNECTED_2522, SV2V_UNCONNECTED_2523, SV2V_UNCONNECTED_2524, SV2V_UNCONNECTED_2525, SV2V_UNCONNECTED_2526, SV2V_UNCONNECTED_2527, SV2V_UNCONNECTED_2528, SV2V_UNCONNECTED_2529, SV2V_UNCONNECTED_2530, SV2V_UNCONNECTED_2531, SV2V_UNCONNECTED_2532, SV2V_UNCONNECTED_2533, SV2V_UNCONNECTED_2534, SV2V_UNCONNECTED_2535, SV2V_UNCONNECTED_2536, SV2V_UNCONNECTED_2537, SV2V_UNCONNECTED_2538, SV2V_UNCONNECTED_2539, SV2V_UNCONNECTED_2540, SV2V_UNCONNECTED_2541, SV2V_UNCONNECTED_2542, SV2V_UNCONNECTED_2543, SV2V_UNCONNECTED_2544, SV2V_UNCONNECTED_2545, SV2V_UNCONNECTED_2546, SV2V_UNCONNECTED_2547, SV2V_UNCONNECTED_2548, SV2V_UNCONNECTED_2549, SV2V_UNCONNECTED_2550, SV2V_UNCONNECTED_2551, SV2V_UNCONNECTED_2552, SV2V_UNCONNECTED_2553, SV2V_UNCONNECTED_2554, SV2V_UNCONNECTED_2555, SV2V_UNCONNECTED_2556, SV2V_UNCONNECTED_2557, SV2V_UNCONNECTED_2558, SV2V_UNCONNECTED_2559, SV2V_UNCONNECTED_2560, SV2V_UNCONNECTED_2561, SV2V_UNCONNECTED_2562, SV2V_UNCONNECTED_2563, SV2V_UNCONNECTED_2564, SV2V_UNCONNECTED_2565, SV2V_UNCONNECTED_2566, SV2V_UNCONNECTED_2567, SV2V_UNCONNECTED_2568, SV2V_UNCONNECTED_2569, SV2V_UNCONNECTED_2570, SV2V_UNCONNECTED_2571, SV2V_UNCONNECTED_2572, SV2V_UNCONNECTED_2573, SV2V_UNCONNECTED_2574, SV2V_UNCONNECTED_2575, SV2V_UNCONNECTED_2576, SV2V_UNCONNECTED_2577, SV2V_UNCONNECTED_2578, SV2V_UNCONNECTED_2579, SV2V_UNCONNECTED_2580, SV2V_UNCONNECTED_2581, SV2V_UNCONNECTED_2582, SV2V_UNCONNECTED_2583, SV2V_UNCONNECTED_2584, SV2V_UNCONNECTED_2585, SV2V_UNCONNECTED_2586, SV2V_UNCONNECTED_2587, SV2V_UNCONNECTED_2588, SV2V_UNCONNECTED_2589, SV2V_UNCONNECTED_2590, SV2V_UNCONNECTED_2591, SV2V_UNCONNECTED_2592, SV2V_UNCONNECTED_2593, SV2V_UNCONNECTED_2594, SV2V_UNCONNECTED_2595, SV2V_UNCONNECTED_2596, SV2V_UNCONNECTED_2597, SV2V_UNCONNECTED_2598, SV2V_UNCONNECTED_2599, SV2V_UNCONNECTED_2600, SV2V_UNCONNECTED_2601, SV2V_UNCONNECTED_2602, SV2V_UNCONNECTED_2603, SV2V_UNCONNECTED_2604, SV2V_UNCONNECTED_2605, SV2V_UNCONNECTED_2606, SV2V_UNCONNECTED_2607, SV2V_UNCONNECTED_2608, SV2V_UNCONNECTED_2609, SV2V_UNCONNECTED_2610, SV2V_UNCONNECTED_2611, SV2V_UNCONNECTED_2612, SV2V_UNCONNECTED_2613, SV2V_UNCONNECTED_2614, SV2V_UNCONNECTED_2615, SV2V_UNCONNECTED_2616, SV2V_UNCONNECTED_2617, SV2V_UNCONNECTED_2618, SV2V_UNCONNECTED_2619, SV2V_UNCONNECTED_2620, SV2V_UNCONNECTED_2621, SV2V_UNCONNECTED_2622, SV2V_UNCONNECTED_2623, SV2V_UNCONNECTED_2624, SV2V_UNCONNECTED_2625, SV2V_UNCONNECTED_2626, SV2V_UNCONNECTED_2627, SV2V_UNCONNECTED_2628, SV2V_UNCONNECTED_2629, SV2V_UNCONNECTED_2630, SV2V_UNCONNECTED_2631, SV2V_UNCONNECTED_2632, SV2V_UNCONNECTED_2633, SV2V_UNCONNECTED_2634, SV2V_UNCONNECTED_2635, SV2V_UNCONNECTED_2636, SV2V_UNCONNECTED_2637, SV2V_UNCONNECTED_2638, SV2V_UNCONNECTED_2639, SV2V_UNCONNECTED_2640, SV2V_UNCONNECTED_2641, SV2V_UNCONNECTED_2642, SV2V_UNCONNECTED_2643, SV2V_UNCONNECTED_2644, SV2V_UNCONNECTED_2645, SV2V_UNCONNECTED_2646, SV2V_UNCONNECTED_2647, SV2V_UNCONNECTED_2648, SV2V_UNCONNECTED_2649, SV2V_UNCONNECTED_2650, SV2V_UNCONNECTED_2651, SV2V_UNCONNECTED_2652, SV2V_UNCONNECTED_2653, SV2V_UNCONNECTED_2654, SV2V_UNCONNECTED_2655, SV2V_UNCONNECTED_2656, SV2V_UNCONNECTED_2657, SV2V_UNCONNECTED_2658, SV2V_UNCONNECTED_2659, SV2V_UNCONNECTED_2660, SV2V_UNCONNECTED_2661, SV2V_UNCONNECTED_2662, SV2V_UNCONNECTED_2663, SV2V_UNCONNECTED_2664, SV2V_UNCONNECTED_2665, SV2V_UNCONNECTED_2666, SV2V_UNCONNECTED_2667, SV2V_UNCONNECTED_2668, SV2V_UNCONNECTED_2669, SV2V_UNCONNECTED_2670, SV2V_UNCONNECTED_2671, SV2V_UNCONNECTED_2672, SV2V_UNCONNECTED_2673, SV2V_UNCONNECTED_2674, SV2V_UNCONNECTED_2675, SV2V_UNCONNECTED_2676, SV2V_UNCONNECTED_2677, SV2V_UNCONNECTED_2678, SV2V_UNCONNECTED_2679, SV2V_UNCONNECTED_2680, SV2V_UNCONNECTED_2681, SV2V_UNCONNECTED_2682, SV2V_UNCONNECTED_2683, SV2V_UNCONNECTED_2684, SV2V_UNCONNECTED_2685, SV2V_UNCONNECTED_2686, SV2V_UNCONNECTED_2687, SV2V_UNCONNECTED_2688, SV2V_UNCONNECTED_2689, SV2V_UNCONNECTED_2690, SV2V_UNCONNECTED_2691, SV2V_UNCONNECTED_2692, SV2V_UNCONNECTED_2693, SV2V_UNCONNECTED_2694, SV2V_UNCONNECTED_2695, SV2V_UNCONNECTED_2696, SV2V_UNCONNECTED_2697, SV2V_UNCONNECTED_2698, SV2V_UNCONNECTED_2699, SV2V_UNCONNECTED_2700, SV2V_UNCONNECTED_2701, SV2V_UNCONNECTED_2702, SV2V_UNCONNECTED_2703, SV2V_UNCONNECTED_2704, SV2V_UNCONNECTED_2705, SV2V_UNCONNECTED_2706, SV2V_UNCONNECTED_2707, SV2V_UNCONNECTED_2708, SV2V_UNCONNECTED_2709, SV2V_UNCONNECTED_2710, SV2V_UNCONNECTED_2711, SV2V_UNCONNECTED_2712, SV2V_UNCONNECTED_2713, SV2V_UNCONNECTED_2714, SV2V_UNCONNECTED_2715, SV2V_UNCONNECTED_2716, SV2V_UNCONNECTED_2717, SV2V_UNCONNECTED_2718, SV2V_UNCONNECTED_2719, SV2V_UNCONNECTED_2720, SV2V_UNCONNECTED_2721, SV2V_UNCONNECTED_2722, SV2V_UNCONNECTED_2723, SV2V_UNCONNECTED_2724, SV2V_UNCONNECTED_2725, SV2V_UNCONNECTED_2726, SV2V_UNCONNECTED_2727, SV2V_UNCONNECTED_2728, SV2V_UNCONNECTED_2729, SV2V_UNCONNECTED_2730, SV2V_UNCONNECTED_2731, SV2V_UNCONNECTED_2732, SV2V_UNCONNECTED_2733, SV2V_UNCONNECTED_2734, SV2V_UNCONNECTED_2735, SV2V_UNCONNECTED_2736, SV2V_UNCONNECTED_2737, SV2V_UNCONNECTED_2738, SV2V_UNCONNECTED_2739, SV2V_UNCONNECTED_2740, SV2V_UNCONNECTED_2741, SV2V_UNCONNECTED_2742, SV2V_UNCONNECTED_2743, SV2V_UNCONNECTED_2744, SV2V_UNCONNECTED_2745, SV2V_UNCONNECTED_2746, SV2V_UNCONNECTED_2747, SV2V_UNCONNECTED_2748, SV2V_UNCONNECTED_2749, SV2V_UNCONNECTED_2750, SV2V_UNCONNECTED_2751, SV2V_UNCONNECTED_2752, SV2V_UNCONNECTED_2753, SV2V_UNCONNECTED_2754, SV2V_UNCONNECTED_2755, SV2V_UNCONNECTED_2756, SV2V_UNCONNECTED_2757, SV2V_UNCONNECTED_2758, SV2V_UNCONNECTED_2759, SV2V_UNCONNECTED_2760, SV2V_UNCONNECTED_2761, SV2V_UNCONNECTED_2762, SV2V_UNCONNECTED_2763, SV2V_UNCONNECTED_2764, SV2V_UNCONNECTED_2765, SV2V_UNCONNECTED_2766, SV2V_UNCONNECTED_2767, SV2V_UNCONNECTED_2768, SV2V_UNCONNECTED_2769, SV2V_UNCONNECTED_2770, SV2V_UNCONNECTED_2771, SV2V_UNCONNECTED_2772, SV2V_UNCONNECTED_2773, SV2V_UNCONNECTED_2774, SV2V_UNCONNECTED_2775, SV2V_UNCONNECTED_2776, SV2V_UNCONNECTED_2777, SV2V_UNCONNECTED_2778, SV2V_UNCONNECTED_2779, SV2V_UNCONNECTED_2780, SV2V_UNCONNECTED_2781, SV2V_UNCONNECTED_2782, SV2V_UNCONNECTED_2783, SV2V_UNCONNECTED_2784, SV2V_UNCONNECTED_2785, SV2V_UNCONNECTED_2786, SV2V_UNCONNECTED_2787, SV2V_UNCONNECTED_2788, SV2V_UNCONNECTED_2789, SV2V_UNCONNECTED_2790, SV2V_UNCONNECTED_2791, SV2V_UNCONNECTED_2792, SV2V_UNCONNECTED_2793, SV2V_UNCONNECTED_2794, SV2V_UNCONNECTED_2795, SV2V_UNCONNECTED_2796, SV2V_UNCONNECTED_2797, SV2V_UNCONNECTED_2798, SV2V_UNCONNECTED_2799, SV2V_UNCONNECTED_2800, SV2V_UNCONNECTED_2801, SV2V_UNCONNECTED_2802, SV2V_UNCONNECTED_2803, SV2V_UNCONNECTED_2804, SV2V_UNCONNECTED_2805, SV2V_UNCONNECTED_2806, SV2V_UNCONNECTED_2807, SV2V_UNCONNECTED_2808, SV2V_UNCONNECTED_2809, SV2V_UNCONNECTED_2810, SV2V_UNCONNECTED_2811, SV2V_UNCONNECTED_2812, SV2V_UNCONNECTED_2813, SV2V_UNCONNECTED_2814, SV2V_UNCONNECTED_2815, SV2V_UNCONNECTED_2816, SV2V_UNCONNECTED_2817, SV2V_UNCONNECTED_2818, SV2V_UNCONNECTED_2819, SV2V_UNCONNECTED_2820, SV2V_UNCONNECTED_2821, SV2V_UNCONNECTED_2822, SV2V_UNCONNECTED_2823, SV2V_UNCONNECTED_2824, SV2V_UNCONNECTED_2825, SV2V_UNCONNECTED_2826, SV2V_UNCONNECTED_2827, SV2V_UNCONNECTED_2828, SV2V_UNCONNECTED_2829, SV2V_UNCONNECTED_2830, SV2V_UNCONNECTED_2831, SV2V_UNCONNECTED_2832, SV2V_UNCONNECTED_2833, SV2V_UNCONNECTED_2834, SV2V_UNCONNECTED_2835, SV2V_UNCONNECTED_2836, SV2V_UNCONNECTED_2837, SV2V_UNCONNECTED_2838, SV2V_UNCONNECTED_2839, SV2V_UNCONNECTED_2840, SV2V_UNCONNECTED_2841, SV2V_UNCONNECTED_2842, SV2V_UNCONNECTED_2843, SV2V_UNCONNECTED_2844, SV2V_UNCONNECTED_2845, SV2V_UNCONNECTED_2846, SV2V_UNCONNECTED_2847, SV2V_UNCONNECTED_2848, SV2V_UNCONNECTED_2849, SV2V_UNCONNECTED_2850, SV2V_UNCONNECTED_2851, SV2V_UNCONNECTED_2852, SV2V_UNCONNECTED_2853, SV2V_UNCONNECTED_2854, SV2V_UNCONNECTED_2855, SV2V_UNCONNECTED_2856, SV2V_UNCONNECTED_2857, SV2V_UNCONNECTED_2858, SV2V_UNCONNECTED_2859, SV2V_UNCONNECTED_2860, SV2V_UNCONNECTED_2861, SV2V_UNCONNECTED_2862, SV2V_UNCONNECTED_2863, SV2V_UNCONNECTED_2864, SV2V_UNCONNECTED_2865, SV2V_UNCONNECTED_2866, SV2V_UNCONNECTED_2867, SV2V_UNCONNECTED_2868, SV2V_UNCONNECTED_2869, SV2V_UNCONNECTED_2870, SV2V_UNCONNECTED_2871, SV2V_UNCONNECTED_2872, SV2V_UNCONNECTED_2873, SV2V_UNCONNECTED_2874, SV2V_UNCONNECTED_2875, SV2V_UNCONNECTED_2876, SV2V_UNCONNECTED_2877, SV2V_UNCONNECTED_2878, SV2V_UNCONNECTED_2879, SV2V_UNCONNECTED_2880, SV2V_UNCONNECTED_2881, SV2V_UNCONNECTED_2882, SV2V_UNCONNECTED_2883, SV2V_UNCONNECTED_2884, SV2V_UNCONNECTED_2885, SV2V_UNCONNECTED_2886, SV2V_UNCONNECTED_2887, SV2V_UNCONNECTED_2888, SV2V_UNCONNECTED_2889, SV2V_UNCONNECTED_2890, SV2V_UNCONNECTED_2891, SV2V_UNCONNECTED_2892, SV2V_UNCONNECTED_2893, SV2V_UNCONNECTED_2894, SV2V_UNCONNECTED_2895, SV2V_UNCONNECTED_2896, SV2V_UNCONNECTED_2897, SV2V_UNCONNECTED_2898, SV2V_UNCONNECTED_2899, SV2V_UNCONNECTED_2900, SV2V_UNCONNECTED_2901, SV2V_UNCONNECTED_2902, SV2V_UNCONNECTED_2903, SV2V_UNCONNECTED_2904, SV2V_UNCONNECTED_2905, SV2V_UNCONNECTED_2906, SV2V_UNCONNECTED_2907, SV2V_UNCONNECTED_2908, SV2V_UNCONNECTED_2909, SV2V_UNCONNECTED_2910, SV2V_UNCONNECTED_2911, SV2V_UNCONNECTED_2912, SV2V_UNCONNECTED_2913, SV2V_UNCONNECTED_2914, SV2V_UNCONNECTED_2915, SV2V_UNCONNECTED_2916, SV2V_UNCONNECTED_2917, SV2V_UNCONNECTED_2918, SV2V_UNCONNECTED_2919, SV2V_UNCONNECTED_2920, SV2V_UNCONNECTED_2921, SV2V_UNCONNECTED_2922, SV2V_UNCONNECTED_2923, SV2V_UNCONNECTED_2924, SV2V_UNCONNECTED_2925, SV2V_UNCONNECTED_2926, SV2V_UNCONNECTED_2927, SV2V_UNCONNECTED_2928, SV2V_UNCONNECTED_2929, SV2V_UNCONNECTED_2930, SV2V_UNCONNECTED_2931, SV2V_UNCONNECTED_2932, SV2V_UNCONNECTED_2933, SV2V_UNCONNECTED_2934, SV2V_UNCONNECTED_2935, SV2V_UNCONNECTED_2936, SV2V_UNCONNECTED_2937, SV2V_UNCONNECTED_2938, SV2V_UNCONNECTED_2939, SV2V_UNCONNECTED_2940, SV2V_UNCONNECTED_2941, SV2V_UNCONNECTED_2942, SV2V_UNCONNECTED_2943, SV2V_UNCONNECTED_2944, SV2V_UNCONNECTED_2945, SV2V_UNCONNECTED_2946, SV2V_UNCONNECTED_2947, SV2V_UNCONNECTED_2948, SV2V_UNCONNECTED_2949, SV2V_UNCONNECTED_2950, SV2V_UNCONNECTED_2951, SV2V_UNCONNECTED_2952, SV2V_UNCONNECTED_2953, SV2V_UNCONNECTED_2954, SV2V_UNCONNECTED_2955, SV2V_UNCONNECTED_2956, SV2V_UNCONNECTED_2957, SV2V_UNCONNECTED_2958, SV2V_UNCONNECTED_2959, SV2V_UNCONNECTED_2960, SV2V_UNCONNECTED_2961, SV2V_UNCONNECTED_2962, SV2V_UNCONNECTED_2963, SV2V_UNCONNECTED_2964, SV2V_UNCONNECTED_2965, SV2V_UNCONNECTED_2966, SV2V_UNCONNECTED_2967, SV2V_UNCONNECTED_2968, SV2V_UNCONNECTED_2969, SV2V_UNCONNECTED_2970, SV2V_UNCONNECTED_2971, SV2V_UNCONNECTED_2972, SV2V_UNCONNECTED_2973, SV2V_UNCONNECTED_2974, SV2V_UNCONNECTED_2975, SV2V_UNCONNECTED_2976, SV2V_UNCONNECTED_2977, SV2V_UNCONNECTED_2978, SV2V_UNCONNECTED_2979, SV2V_UNCONNECTED_2980, SV2V_UNCONNECTED_2981, SV2V_UNCONNECTED_2982, SV2V_UNCONNECTED_2983, SV2V_UNCONNECTED_2984, SV2V_UNCONNECTED_2985, SV2V_UNCONNECTED_2986, SV2V_UNCONNECTED_2987, SV2V_UNCONNECTED_2988, SV2V_UNCONNECTED_2989, SV2V_UNCONNECTED_2990, SV2V_UNCONNECTED_2991, SV2V_UNCONNECTED_2992, SV2V_UNCONNECTED_2993, SV2V_UNCONNECTED_2994, SV2V_UNCONNECTED_2995, SV2V_UNCONNECTED_2996, SV2V_UNCONNECTED_2997, SV2V_UNCONNECTED_2998, SV2V_UNCONNECTED_2999, SV2V_UNCONNECTED_3000, SV2V_UNCONNECTED_3001, SV2V_UNCONNECTED_3002, SV2V_UNCONNECTED_3003, SV2V_UNCONNECTED_3004, SV2V_UNCONNECTED_3005, SV2V_UNCONNECTED_3006, SV2V_UNCONNECTED_3007, SV2V_UNCONNECTED_3008, SV2V_UNCONNECTED_3009, SV2V_UNCONNECTED_3010, SV2V_UNCONNECTED_3011, SV2V_UNCONNECTED_3012, SV2V_UNCONNECTED_3013, SV2V_UNCONNECTED_3014, SV2V_UNCONNECTED_3015, SV2V_UNCONNECTED_3016, SV2V_UNCONNECTED_3017, SV2V_UNCONNECTED_3018, SV2V_UNCONNECTED_3019, SV2V_UNCONNECTED_3020, SV2V_UNCONNECTED_3021, SV2V_UNCONNECTED_3022, SV2V_UNCONNECTED_3023, SV2V_UNCONNECTED_3024, SV2V_UNCONNECTED_3025, SV2V_UNCONNECTED_3026, SV2V_UNCONNECTED_3027, SV2V_UNCONNECTED_3028, SV2V_UNCONNECTED_3029, SV2V_UNCONNECTED_3030, SV2V_UNCONNECTED_3031, SV2V_UNCONNECTED_3032, SV2V_UNCONNECTED_3033, SV2V_UNCONNECTED_3034, SV2V_UNCONNECTED_3035, SV2V_UNCONNECTED_3036, SV2V_UNCONNECTED_3037, SV2V_UNCONNECTED_3038, SV2V_UNCONNECTED_3039, SV2V_UNCONNECTED_3040, SV2V_UNCONNECTED_3041, SV2V_UNCONNECTED_3042, SV2V_UNCONNECTED_3043, SV2V_UNCONNECTED_3044, SV2V_UNCONNECTED_3045, SV2V_UNCONNECTED_3046, SV2V_UNCONNECTED_3047, SV2V_UNCONNECTED_3048, SV2V_UNCONNECTED_3049, SV2V_UNCONNECTED_3050, SV2V_UNCONNECTED_3051, SV2V_UNCONNECTED_3052, SV2V_UNCONNECTED_3053, SV2V_UNCONNECTED_3054, SV2V_UNCONNECTED_3055, SV2V_UNCONNECTED_3056, SV2V_UNCONNECTED_3057, SV2V_UNCONNECTED_3058, SV2V_UNCONNECTED_3059, SV2V_UNCONNECTED_3060, SV2V_UNCONNECTED_3061, SV2V_UNCONNECTED_3062, SV2V_UNCONNECTED_3063, SV2V_UNCONNECTED_3064, SV2V_UNCONNECTED_3065, SV2V_UNCONNECTED_3066, SV2V_UNCONNECTED_3067, SV2V_UNCONNECTED_3068, SV2V_UNCONNECTED_3069, SV2V_UNCONNECTED_3070, SV2V_UNCONNECTED_3071, SV2V_UNCONNECTED_3072, SV2V_UNCONNECTED_3073, SV2V_UNCONNECTED_3074, SV2V_UNCONNECTED_3075, SV2V_UNCONNECTED_3076, SV2V_UNCONNECTED_3077, SV2V_UNCONNECTED_3078, SV2V_UNCONNECTED_3079, SV2V_UNCONNECTED_3080, SV2V_UNCONNECTED_3081, SV2V_UNCONNECTED_3082, SV2V_UNCONNECTED_3083, SV2V_UNCONNECTED_3084, SV2V_UNCONNECTED_3085, SV2V_UNCONNECTED_3086, SV2V_UNCONNECTED_3087, SV2V_UNCONNECTED_3088, SV2V_UNCONNECTED_3089, SV2V_UNCONNECTED_3090, SV2V_UNCONNECTED_3091, SV2V_UNCONNECTED_3092, SV2V_UNCONNECTED_3093, SV2V_UNCONNECTED_3094, SV2V_UNCONNECTED_3095, SV2V_UNCONNECTED_3096, SV2V_UNCONNECTED_3097, SV2V_UNCONNECTED_3098, SV2V_UNCONNECTED_3099, SV2V_UNCONNECTED_3100, SV2V_UNCONNECTED_3101, SV2V_UNCONNECTED_3102, SV2V_UNCONNECTED_3103, SV2V_UNCONNECTED_3104, SV2V_UNCONNECTED_3105, SV2V_UNCONNECTED_3106, SV2V_UNCONNECTED_3107, SV2V_UNCONNECTED_3108, SV2V_UNCONNECTED_3109, SV2V_UNCONNECTED_3110, SV2V_UNCONNECTED_3111, SV2V_UNCONNECTED_3112, SV2V_UNCONNECTED_3113, SV2V_UNCONNECTED_3114, SV2V_UNCONNECTED_3115, SV2V_UNCONNECTED_3116, SV2V_UNCONNECTED_3117, SV2V_UNCONNECTED_3118, SV2V_UNCONNECTED_3119, SV2V_UNCONNECTED_3120, SV2V_UNCONNECTED_3121, SV2V_UNCONNECTED_3122, SV2V_UNCONNECTED_3123, SV2V_UNCONNECTED_3124, SV2V_UNCONNECTED_3125, SV2V_UNCONNECTED_3126, SV2V_UNCONNECTED_3127, SV2V_UNCONNECTED_3128, SV2V_UNCONNECTED_3129, SV2V_UNCONNECTED_3130, SV2V_UNCONNECTED_3131, SV2V_UNCONNECTED_3132, SV2V_UNCONNECTED_3133, SV2V_UNCONNECTED_3134, SV2V_UNCONNECTED_3135, SV2V_UNCONNECTED_3136, SV2V_UNCONNECTED_3137, SV2V_UNCONNECTED_3138, SV2V_UNCONNECTED_3139, SV2V_UNCONNECTED_3140, SV2V_UNCONNECTED_3141, SV2V_UNCONNECTED_3142, SV2V_UNCONNECTED_3143, SV2V_UNCONNECTED_3144, SV2V_UNCONNECTED_3145, SV2V_UNCONNECTED_3146, SV2V_UNCONNECTED_3147, SV2V_UNCONNECTED_3148, SV2V_UNCONNECTED_3149, SV2V_UNCONNECTED_3150, SV2V_UNCONNECTED_3151, SV2V_UNCONNECTED_3152, SV2V_UNCONNECTED_3153, SV2V_UNCONNECTED_3154, SV2V_UNCONNECTED_3155, SV2V_UNCONNECTED_3156, SV2V_UNCONNECTED_3157, SV2V_UNCONNECTED_3158, SV2V_UNCONNECTED_3159, SV2V_UNCONNECTED_3160, SV2V_UNCONNECTED_3161, SV2V_UNCONNECTED_3162, SV2V_UNCONNECTED_3163, SV2V_UNCONNECTED_3164, SV2V_UNCONNECTED_3165, SV2V_UNCONNECTED_3166, SV2V_UNCONNECTED_3167, SV2V_UNCONNECTED_3168, SV2V_UNCONNECTED_3169, SV2V_UNCONNECTED_3170, SV2V_UNCONNECTED_3171, SV2V_UNCONNECTED_3172, SV2V_UNCONNECTED_3173, SV2V_UNCONNECTED_3174, SV2V_UNCONNECTED_3175, SV2V_UNCONNECTED_3176, SV2V_UNCONNECTED_3177, SV2V_UNCONNECTED_3178, SV2V_UNCONNECTED_3179, SV2V_UNCONNECTED_3180, SV2V_UNCONNECTED_3181, SV2V_UNCONNECTED_3182, SV2V_UNCONNECTED_3183, SV2V_UNCONNECTED_3184, SV2V_UNCONNECTED_3185, SV2V_UNCONNECTED_3186, SV2V_UNCONNECTED_3187, SV2V_UNCONNECTED_3188, SV2V_UNCONNECTED_3189, SV2V_UNCONNECTED_3190, SV2V_UNCONNECTED_3191, SV2V_UNCONNECTED_3192, SV2V_UNCONNECTED_3193, SV2V_UNCONNECTED_3194, SV2V_UNCONNECTED_3195, SV2V_UNCONNECTED_3196, SV2V_UNCONNECTED_3197, SV2V_UNCONNECTED_3198, SV2V_UNCONNECTED_3199, SV2V_UNCONNECTED_3200, SV2V_UNCONNECTED_3201, SV2V_UNCONNECTED_3202, SV2V_UNCONNECTED_3203, SV2V_UNCONNECTED_3204, SV2V_UNCONNECTED_3205, SV2V_UNCONNECTED_3206, SV2V_UNCONNECTED_3207, SV2V_UNCONNECTED_3208, SV2V_UNCONNECTED_3209, SV2V_UNCONNECTED_3210, SV2V_UNCONNECTED_3211, SV2V_UNCONNECTED_3212, SV2V_UNCONNECTED_3213, SV2V_UNCONNECTED_3214, SV2V_UNCONNECTED_3215, SV2V_UNCONNECTED_3216, SV2V_UNCONNECTED_3217, SV2V_UNCONNECTED_3218, SV2V_UNCONNECTED_3219, SV2V_UNCONNECTED_3220, SV2V_UNCONNECTED_3221, SV2V_UNCONNECTED_3222, SV2V_UNCONNECTED_3223, SV2V_UNCONNECTED_3224, SV2V_UNCONNECTED_3225, SV2V_UNCONNECTED_3226, SV2V_UNCONNECTED_3227, SV2V_UNCONNECTED_3228, SV2V_UNCONNECTED_3229, SV2V_UNCONNECTED_3230, SV2V_UNCONNECTED_3231, SV2V_UNCONNECTED_3232, SV2V_UNCONNECTED_3233, SV2V_UNCONNECTED_3234, SV2V_UNCONNECTED_3235, SV2V_UNCONNECTED_3236, SV2V_UNCONNECTED_3237, SV2V_UNCONNECTED_3238, SV2V_UNCONNECTED_3239, SV2V_UNCONNECTED_3240, SV2V_UNCONNECTED_3241, SV2V_UNCONNECTED_3242, SV2V_UNCONNECTED_3243, SV2V_UNCONNECTED_3244, SV2V_UNCONNECTED_3245, SV2V_UNCONNECTED_3246, SV2V_UNCONNECTED_3247, SV2V_UNCONNECTED_3248, SV2V_UNCONNECTED_3249, SV2V_UNCONNECTED_3250, SV2V_UNCONNECTED_3251, SV2V_UNCONNECTED_3252, SV2V_UNCONNECTED_3253, SV2V_UNCONNECTED_3254, SV2V_UNCONNECTED_3255, SV2V_UNCONNECTED_3256, SV2V_UNCONNECTED_3257, SV2V_UNCONNECTED_3258, SV2V_UNCONNECTED_3259, SV2V_UNCONNECTED_3260, SV2V_UNCONNECTED_3261, SV2V_UNCONNECTED_3262, SV2V_UNCONNECTED_3263, SV2V_UNCONNECTED_3264, SV2V_UNCONNECTED_3265, SV2V_UNCONNECTED_3266, SV2V_UNCONNECTED_3267, SV2V_UNCONNECTED_3268, SV2V_UNCONNECTED_3269, SV2V_UNCONNECTED_3270, SV2V_UNCONNECTED_3271, SV2V_UNCONNECTED_3272, SV2V_UNCONNECTED_3273, SV2V_UNCONNECTED_3274, SV2V_UNCONNECTED_3275, SV2V_UNCONNECTED_3276, SV2V_UNCONNECTED_3277, SV2V_UNCONNECTED_3278, SV2V_UNCONNECTED_3279, SV2V_UNCONNECTED_3280, SV2V_UNCONNECTED_3281, SV2V_UNCONNECTED_3282, SV2V_UNCONNECTED_3283, SV2V_UNCONNECTED_3284, SV2V_UNCONNECTED_3285, SV2V_UNCONNECTED_3286, SV2V_UNCONNECTED_3287, SV2V_UNCONNECTED_3288, SV2V_UNCONNECTED_3289, SV2V_UNCONNECTED_3290, SV2V_UNCONNECTED_3291, SV2V_UNCONNECTED_3292, SV2V_UNCONNECTED_3293, SV2V_UNCONNECTED_3294, SV2V_UNCONNECTED_3295, SV2V_UNCONNECTED_3296, SV2V_UNCONNECTED_3297, SV2V_UNCONNECTED_3298, SV2V_UNCONNECTED_3299, SV2V_UNCONNECTED_3300, SV2V_UNCONNECTED_3301, SV2V_UNCONNECTED_3302, SV2V_UNCONNECTED_3303, SV2V_UNCONNECTED_3304, SV2V_UNCONNECTED_3305, SV2V_UNCONNECTED_3306, SV2V_UNCONNECTED_3307, SV2V_UNCONNECTED_3308, SV2V_UNCONNECTED_3309, SV2V_UNCONNECTED_3310, SV2V_UNCONNECTED_3311, SV2V_UNCONNECTED_3312, SV2V_UNCONNECTED_3313, SV2V_UNCONNECTED_3314, SV2V_UNCONNECTED_3315, SV2V_UNCONNECTED_3316, SV2V_UNCONNECTED_3317, SV2V_UNCONNECTED_3318, SV2V_UNCONNECTED_3319, SV2V_UNCONNECTED_3320, SV2V_UNCONNECTED_3321, SV2V_UNCONNECTED_3322, SV2V_UNCONNECTED_3323, SV2V_UNCONNECTED_3324, SV2V_UNCONNECTED_3325, SV2V_UNCONNECTED_3326, SV2V_UNCONNECTED_3327, SV2V_UNCONNECTED_3328, SV2V_UNCONNECTED_3329, SV2V_UNCONNECTED_3330, SV2V_UNCONNECTED_3331, SV2V_UNCONNECTED_3332, SV2V_UNCONNECTED_3333, SV2V_UNCONNECTED_3334, SV2V_UNCONNECTED_3335, SV2V_UNCONNECTED_3336, SV2V_UNCONNECTED_3337, SV2V_UNCONNECTED_3338, SV2V_UNCONNECTED_3339, SV2V_UNCONNECTED_3340, SV2V_UNCONNECTED_3341, SV2V_UNCONNECTED_3342, SV2V_UNCONNECTED_3343, SV2V_UNCONNECTED_3344, SV2V_UNCONNECTED_3345, SV2V_UNCONNECTED_3346, SV2V_UNCONNECTED_3347, SV2V_UNCONNECTED_3348, SV2V_UNCONNECTED_3349, SV2V_UNCONNECTED_3350, SV2V_UNCONNECTED_3351, SV2V_UNCONNECTED_3352, SV2V_UNCONNECTED_3353, SV2V_UNCONNECTED_3354, SV2V_UNCONNECTED_3355, SV2V_UNCONNECTED_3356, SV2V_UNCONNECTED_3357, SV2V_UNCONNECTED_3358, SV2V_UNCONNECTED_3359, SV2V_UNCONNECTED_3360, SV2V_UNCONNECTED_3361, SV2V_UNCONNECTED_3362, SV2V_UNCONNECTED_3363, SV2V_UNCONNECTED_3364, SV2V_UNCONNECTED_3365, SV2V_UNCONNECTED_3366, SV2V_UNCONNECTED_3367, SV2V_UNCONNECTED_3368, SV2V_UNCONNECTED_3369, SV2V_UNCONNECTED_3370, SV2V_UNCONNECTED_3371, SV2V_UNCONNECTED_3372, SV2V_UNCONNECTED_3373, SV2V_UNCONNECTED_3374, SV2V_UNCONNECTED_3375, SV2V_UNCONNECTED_3376, SV2V_UNCONNECTED_3377, SV2V_UNCONNECTED_3378, SV2V_UNCONNECTED_3379, SV2V_UNCONNECTED_3380, SV2V_UNCONNECTED_3381, SV2V_UNCONNECTED_3382, SV2V_UNCONNECTED_3383, SV2V_UNCONNECTED_3384, SV2V_UNCONNECTED_3385, SV2V_UNCONNECTED_3386, SV2V_UNCONNECTED_3387, SV2V_UNCONNECTED_3388, SV2V_UNCONNECTED_3389, SV2V_UNCONNECTED_3390, SV2V_UNCONNECTED_3391, SV2V_UNCONNECTED_3392, SV2V_UNCONNECTED_3393, SV2V_UNCONNECTED_3394, SV2V_UNCONNECTED_3395, SV2V_UNCONNECTED_3396, SV2V_UNCONNECTED_3397, SV2V_UNCONNECTED_3398, SV2V_UNCONNECTED_3399, SV2V_UNCONNECTED_3400, SV2V_UNCONNECTED_3401, SV2V_UNCONNECTED_3402, SV2V_UNCONNECTED_3403, SV2V_UNCONNECTED_3404, SV2V_UNCONNECTED_3405, SV2V_UNCONNECTED_3406, SV2V_UNCONNECTED_3407, SV2V_UNCONNECTED_3408, SV2V_UNCONNECTED_3409, SV2V_UNCONNECTED_3410, SV2V_UNCONNECTED_3411, SV2V_UNCONNECTED_3412, SV2V_UNCONNECTED_3413, SV2V_UNCONNECTED_3414, SV2V_UNCONNECTED_3415, SV2V_UNCONNECTED_3416, SV2V_UNCONNECTED_3417, SV2V_UNCONNECTED_3418, SV2V_UNCONNECTED_3419, SV2V_UNCONNECTED_3420, SV2V_UNCONNECTED_3421, SV2V_UNCONNECTED_3422, SV2V_UNCONNECTED_3423, SV2V_UNCONNECTED_3424, SV2V_UNCONNECTED_3425, SV2V_UNCONNECTED_3426, SV2V_UNCONNECTED_3427, SV2V_UNCONNECTED_3428, SV2V_UNCONNECTED_3429, SV2V_UNCONNECTED_3430, SV2V_UNCONNECTED_3431, SV2V_UNCONNECTED_3432, SV2V_UNCONNECTED_3433, SV2V_UNCONNECTED_3434, SV2V_UNCONNECTED_3435, SV2V_UNCONNECTED_3436, SV2V_UNCONNECTED_3437, SV2V_UNCONNECTED_3438, SV2V_UNCONNECTED_3439, SV2V_UNCONNECTED_3440, SV2V_UNCONNECTED_3441, SV2V_UNCONNECTED_3442, SV2V_UNCONNECTED_3443, SV2V_UNCONNECTED_3444, SV2V_UNCONNECTED_3445, SV2V_UNCONNECTED_3446, SV2V_UNCONNECTED_3447, SV2V_UNCONNECTED_3448, SV2V_UNCONNECTED_3449, SV2V_UNCONNECTED_3450, SV2V_UNCONNECTED_3451, SV2V_UNCONNECTED_3452, SV2V_UNCONNECTED_3453, SV2V_UNCONNECTED_3454, SV2V_UNCONNECTED_3455, SV2V_UNCONNECTED_3456, SV2V_UNCONNECTED_3457, SV2V_UNCONNECTED_3458, SV2V_UNCONNECTED_3459, SV2V_UNCONNECTED_3460, SV2V_UNCONNECTED_3461, SV2V_UNCONNECTED_3462, SV2V_UNCONNECTED_3463, SV2V_UNCONNECTED_3464, SV2V_UNCONNECTED_3465, SV2V_UNCONNECTED_3466, SV2V_UNCONNECTED_3467, SV2V_UNCONNECTED_3468, SV2V_UNCONNECTED_3469, SV2V_UNCONNECTED_3470, SV2V_UNCONNECTED_3471, SV2V_UNCONNECTED_3472, SV2V_UNCONNECTED_3473, SV2V_UNCONNECTED_3474, SV2V_UNCONNECTED_3475, SV2V_UNCONNECTED_3476, SV2V_UNCONNECTED_3477, SV2V_UNCONNECTED_3478, SV2V_UNCONNECTED_3479, SV2V_UNCONNECTED_3480, SV2V_UNCONNECTED_3481, SV2V_UNCONNECTED_3482, SV2V_UNCONNECTED_3483, SV2V_UNCONNECTED_3484, SV2V_UNCONNECTED_3485, SV2V_UNCONNECTED_3486, SV2V_UNCONNECTED_3487, SV2V_UNCONNECTED_3488, SV2V_UNCONNECTED_3489, SV2V_UNCONNECTED_3490, SV2V_UNCONNECTED_3491, SV2V_UNCONNECTED_3492, SV2V_UNCONNECTED_3493, SV2V_UNCONNECTED_3494, SV2V_UNCONNECTED_3495, SV2V_UNCONNECTED_3496, SV2V_UNCONNECTED_3497, SV2V_UNCONNECTED_3498, SV2V_UNCONNECTED_3499, SV2V_UNCONNECTED_3500, SV2V_UNCONNECTED_3501, SV2V_UNCONNECTED_3502, SV2V_UNCONNECTED_3503, SV2V_UNCONNECTED_3504, SV2V_UNCONNECTED_3505, SV2V_UNCONNECTED_3506, SV2V_UNCONNECTED_3507, SV2V_UNCONNECTED_3508, SV2V_UNCONNECTED_3509, SV2V_UNCONNECTED_3510, SV2V_UNCONNECTED_3511, SV2V_UNCONNECTED_3512, SV2V_UNCONNECTED_3513, SV2V_UNCONNECTED_3514, SV2V_UNCONNECTED_3515, SV2V_UNCONNECTED_3516, SV2V_UNCONNECTED_3517, SV2V_UNCONNECTED_3518, SV2V_UNCONNECTED_3519, SV2V_UNCONNECTED_3520, SV2V_UNCONNECTED_3521, SV2V_UNCONNECTED_3522, SV2V_UNCONNECTED_3523, SV2V_UNCONNECTED_3524, SV2V_UNCONNECTED_3525, SV2V_UNCONNECTED_3526, SV2V_UNCONNECTED_3527, SV2V_UNCONNECTED_3528, SV2V_UNCONNECTED_3529, SV2V_UNCONNECTED_3530, SV2V_UNCONNECTED_3531, SV2V_UNCONNECTED_3532, SV2V_UNCONNECTED_3533, SV2V_UNCONNECTED_3534, SV2V_UNCONNECTED_3535, SV2V_UNCONNECTED_3536, SV2V_UNCONNECTED_3537, SV2V_UNCONNECTED_3538, SV2V_UNCONNECTED_3539, SV2V_UNCONNECTED_3540, SV2V_UNCONNECTED_3541, SV2V_UNCONNECTED_3542, SV2V_UNCONNECTED_3543, SV2V_UNCONNECTED_3544, SV2V_UNCONNECTED_3545, SV2V_UNCONNECTED_3546, SV2V_UNCONNECTED_3547, SV2V_UNCONNECTED_3548, SV2V_UNCONNECTED_3549, SV2V_UNCONNECTED_3550, SV2V_UNCONNECTED_3551, SV2V_UNCONNECTED_3552, SV2V_UNCONNECTED_3553, SV2V_UNCONNECTED_3554, SV2V_UNCONNECTED_3555, SV2V_UNCONNECTED_3556, SV2V_UNCONNECTED_3557, SV2V_UNCONNECTED_3558, SV2V_UNCONNECTED_3559, SV2V_UNCONNECTED_3560, SV2V_UNCONNECTED_3561, SV2V_UNCONNECTED_3562, SV2V_UNCONNECTED_3563, SV2V_UNCONNECTED_3564, SV2V_UNCONNECTED_3565, SV2V_UNCONNECTED_3566, SV2V_UNCONNECTED_3567, SV2V_UNCONNECTED_3568, SV2V_UNCONNECTED_3569, SV2V_UNCONNECTED_3570, SV2V_UNCONNECTED_3571, SV2V_UNCONNECTED_3572, SV2V_UNCONNECTED_3573, SV2V_UNCONNECTED_3574, SV2V_UNCONNECTED_3575, SV2V_UNCONNECTED_3576, SV2V_UNCONNECTED_3577, SV2V_UNCONNECTED_3578, SV2V_UNCONNECTED_3579, SV2V_UNCONNECTED_3580, SV2V_UNCONNECTED_3581, SV2V_UNCONNECTED_3582, SV2V_UNCONNECTED_3583, SV2V_UNCONNECTED_3584, SV2V_UNCONNECTED_3585, SV2V_UNCONNECTED_3586, SV2V_UNCONNECTED_3587, SV2V_UNCONNECTED_3588, SV2V_UNCONNECTED_3589, SV2V_UNCONNECTED_3590, SV2V_UNCONNECTED_3591, SV2V_UNCONNECTED_3592, SV2V_UNCONNECTED_3593, SV2V_UNCONNECTED_3594, SV2V_UNCONNECTED_3595, SV2V_UNCONNECTED_3596, SV2V_UNCONNECTED_3597, SV2V_UNCONNECTED_3598, SV2V_UNCONNECTED_3599, SV2V_UNCONNECTED_3600, SV2V_UNCONNECTED_3601, SV2V_UNCONNECTED_3602, SV2V_UNCONNECTED_3603, SV2V_UNCONNECTED_3604, SV2V_UNCONNECTED_3605, SV2V_UNCONNECTED_3606, SV2V_UNCONNECTED_3607, SV2V_UNCONNECTED_3608, SV2V_UNCONNECTED_3609, SV2V_UNCONNECTED_3610, SV2V_UNCONNECTED_3611, SV2V_UNCONNECTED_3612, SV2V_UNCONNECTED_3613, SV2V_UNCONNECTED_3614, SV2V_UNCONNECTED_3615, SV2V_UNCONNECTED_3616, SV2V_UNCONNECTED_3617, SV2V_UNCONNECTED_3618, SV2V_UNCONNECTED_3619, SV2V_UNCONNECTED_3620, SV2V_UNCONNECTED_3621, SV2V_UNCONNECTED_3622, SV2V_UNCONNECTED_3623, SV2V_UNCONNECTED_3624, SV2V_UNCONNECTED_3625, SV2V_UNCONNECTED_3626, SV2V_UNCONNECTED_3627, SV2V_UNCONNECTED_3628, SV2V_UNCONNECTED_3629, SV2V_UNCONNECTED_3630, SV2V_UNCONNECTED_3631, SV2V_UNCONNECTED_3632, SV2V_UNCONNECTED_3633, SV2V_UNCONNECTED_3634, SV2V_UNCONNECTED_3635, SV2V_UNCONNECTED_3636, SV2V_UNCONNECTED_3637, SV2V_UNCONNECTED_3638, SV2V_UNCONNECTED_3639, SV2V_UNCONNECTED_3640, SV2V_UNCONNECTED_3641, SV2V_UNCONNECTED_3642, SV2V_UNCONNECTED_3643, SV2V_UNCONNECTED_3644, SV2V_UNCONNECTED_3645, SV2V_UNCONNECTED_3646, SV2V_UNCONNECTED_3647, SV2V_UNCONNECTED_3648, SV2V_UNCONNECTED_3649, SV2V_UNCONNECTED_3650, SV2V_UNCONNECTED_3651, SV2V_UNCONNECTED_3652, SV2V_UNCONNECTED_3653, SV2V_UNCONNECTED_3654, SV2V_UNCONNECTED_3655, SV2V_UNCONNECTED_3656, SV2V_UNCONNECTED_3657, SV2V_UNCONNECTED_3658, SV2V_UNCONNECTED_3659, SV2V_UNCONNECTED_3660, SV2V_UNCONNECTED_3661, SV2V_UNCONNECTED_3662, SV2V_UNCONNECTED_3663, SV2V_UNCONNECTED_3664, SV2V_UNCONNECTED_3665, SV2V_UNCONNECTED_3666, SV2V_UNCONNECTED_3667, SV2V_UNCONNECTED_3668, SV2V_UNCONNECTED_3669, SV2V_UNCONNECTED_3670, SV2V_UNCONNECTED_3671, SV2V_UNCONNECTED_3672, SV2V_UNCONNECTED_3673, SV2V_UNCONNECTED_3674, SV2V_UNCONNECTED_3675, SV2V_UNCONNECTED_3676, SV2V_UNCONNECTED_3677, SV2V_UNCONNECTED_3678, SV2V_UNCONNECTED_3679, SV2V_UNCONNECTED_3680, SV2V_UNCONNECTED_3681, SV2V_UNCONNECTED_3682, SV2V_UNCONNECTED_3683, SV2V_UNCONNECTED_3684, SV2V_UNCONNECTED_3685, SV2V_UNCONNECTED_3686, SV2V_UNCONNECTED_3687, SV2V_UNCONNECTED_3688, SV2V_UNCONNECTED_3689, SV2V_UNCONNECTED_3690, SV2V_UNCONNECTED_3691, SV2V_UNCONNECTED_3692, SV2V_UNCONNECTED_3693, SV2V_UNCONNECTED_3694, SV2V_UNCONNECTED_3695, SV2V_UNCONNECTED_3696, SV2V_UNCONNECTED_3697, SV2V_UNCONNECTED_3698, SV2V_UNCONNECTED_3699, SV2V_UNCONNECTED_3700, SV2V_UNCONNECTED_3701, SV2V_UNCONNECTED_3702, SV2V_UNCONNECTED_3703, SV2V_UNCONNECTED_3704, SV2V_UNCONNECTED_3705, SV2V_UNCONNECTED_3706, SV2V_UNCONNECTED_3707, SV2V_UNCONNECTED_3708, SV2V_UNCONNECTED_3709, SV2V_UNCONNECTED_3710, SV2V_UNCONNECTED_3711, SV2V_UNCONNECTED_3712, SV2V_UNCONNECTED_3713, SV2V_UNCONNECTED_3714, SV2V_UNCONNECTED_3715, SV2V_UNCONNECTED_3716, SV2V_UNCONNECTED_3717, SV2V_UNCONNECTED_3718, SV2V_UNCONNECTED_3719, SV2V_UNCONNECTED_3720, SV2V_UNCONNECTED_3721, SV2V_UNCONNECTED_3722, SV2V_UNCONNECTED_3723, SV2V_UNCONNECTED_3724, SV2V_UNCONNECTED_3725, SV2V_UNCONNECTED_3726, SV2V_UNCONNECTED_3727, SV2V_UNCONNECTED_3728, SV2V_UNCONNECTED_3729, SV2V_UNCONNECTED_3730, SV2V_UNCONNECTED_3731, SV2V_UNCONNECTED_3732, SV2V_UNCONNECTED_3733, SV2V_UNCONNECTED_3734, SV2V_UNCONNECTED_3735, SV2V_UNCONNECTED_3736, SV2V_UNCONNECTED_3737, SV2V_UNCONNECTED_3738, SV2V_UNCONNECTED_3739, SV2V_UNCONNECTED_3740, SV2V_UNCONNECTED_3741, SV2V_UNCONNECTED_3742, SV2V_UNCONNECTED_3743, SV2V_UNCONNECTED_3744, SV2V_UNCONNECTED_3745, SV2V_UNCONNECTED_3746, SV2V_UNCONNECTED_3747, SV2V_UNCONNECTED_3748, SV2V_UNCONNECTED_3749, SV2V_UNCONNECTED_3750, SV2V_UNCONNECTED_3751, SV2V_UNCONNECTED_3752, SV2V_UNCONNECTED_3753, SV2V_UNCONNECTED_3754, SV2V_UNCONNECTED_3755, SV2V_UNCONNECTED_3756, SV2V_UNCONNECTED_3757, SV2V_UNCONNECTED_3758, SV2V_UNCONNECTED_3759, SV2V_UNCONNECTED_3760, SV2V_UNCONNECTED_3761, SV2V_UNCONNECTED_3762, SV2V_UNCONNECTED_3763, SV2V_UNCONNECTED_3764, SV2V_UNCONNECTED_3765, SV2V_UNCONNECTED_3766, SV2V_UNCONNECTED_3767, SV2V_UNCONNECTED_3768, SV2V_UNCONNECTED_3769, SV2V_UNCONNECTED_3770, SV2V_UNCONNECTED_3771, SV2V_UNCONNECTED_3772, SV2V_UNCONNECTED_3773, SV2V_UNCONNECTED_3774, SV2V_UNCONNECTED_3775, SV2V_UNCONNECTED_3776, SV2V_UNCONNECTED_3777, SV2V_UNCONNECTED_3778, SV2V_UNCONNECTED_3779, SV2V_UNCONNECTED_3780, SV2V_UNCONNECTED_3781, SV2V_UNCONNECTED_3782, SV2V_UNCONNECTED_3783, SV2V_UNCONNECTED_3784, SV2V_UNCONNECTED_3785, SV2V_UNCONNECTED_3786, SV2V_UNCONNECTED_3787, SV2V_UNCONNECTED_3788, SV2V_UNCONNECTED_3789, SV2V_UNCONNECTED_3790, SV2V_UNCONNECTED_3791, SV2V_UNCONNECTED_3792, SV2V_UNCONNECTED_3793, SV2V_UNCONNECTED_3794, SV2V_UNCONNECTED_3795, SV2V_UNCONNECTED_3796, SV2V_UNCONNECTED_3797, SV2V_UNCONNECTED_3798, SV2V_UNCONNECTED_3799, SV2V_UNCONNECTED_3800, SV2V_UNCONNECTED_3801, SV2V_UNCONNECTED_3802, SV2V_UNCONNECTED_3803, SV2V_UNCONNECTED_3804, SV2V_UNCONNECTED_3805, SV2V_UNCONNECTED_3806, SV2V_UNCONNECTED_3807, SV2V_UNCONNECTED_3808, SV2V_UNCONNECTED_3809, SV2V_UNCONNECTED_3810, SV2V_UNCONNECTED_3811, SV2V_UNCONNECTED_3812, SV2V_UNCONNECTED_3813, SV2V_UNCONNECTED_3814, SV2V_UNCONNECTED_3815, SV2V_UNCONNECTED_3816, SV2V_UNCONNECTED_3817, SV2V_UNCONNECTED_3818, SV2V_UNCONNECTED_3819, SV2V_UNCONNECTED_3820, SV2V_UNCONNECTED_3821, SV2V_UNCONNECTED_3822, SV2V_UNCONNECTED_3823, SV2V_UNCONNECTED_3824, SV2V_UNCONNECTED_3825, SV2V_UNCONNECTED_3826, SV2V_UNCONNECTED_3827, SV2V_UNCONNECTED_3828, SV2V_UNCONNECTED_3829, SV2V_UNCONNECTED_3830, SV2V_UNCONNECTED_3831, SV2V_UNCONNECTED_3832, SV2V_UNCONNECTED_3833, SV2V_UNCONNECTED_3834, SV2V_UNCONNECTED_3835, SV2V_UNCONNECTED_3836, SV2V_UNCONNECTED_3837, SV2V_UNCONNECTED_3838, SV2V_UNCONNECTED_3839, SV2V_UNCONNECTED_3840, SV2V_UNCONNECTED_3841, SV2V_UNCONNECTED_3842, SV2V_UNCONNECTED_3843, SV2V_UNCONNECTED_3844, SV2V_UNCONNECTED_3845, SV2V_UNCONNECTED_3846, SV2V_UNCONNECTED_3847, SV2V_UNCONNECTED_3848, SV2V_UNCONNECTED_3849, SV2V_UNCONNECTED_3850, SV2V_UNCONNECTED_3851, SV2V_UNCONNECTED_3852, SV2V_UNCONNECTED_3853, SV2V_UNCONNECTED_3854, SV2V_UNCONNECTED_3855, SV2V_UNCONNECTED_3856, SV2V_UNCONNECTED_3857, SV2V_UNCONNECTED_3858, SV2V_UNCONNECTED_3859, SV2V_UNCONNECTED_3860, SV2V_UNCONNECTED_3861, SV2V_UNCONNECTED_3862, SV2V_UNCONNECTED_3863, SV2V_UNCONNECTED_3864, SV2V_UNCONNECTED_3865, SV2V_UNCONNECTED_3866, SV2V_UNCONNECTED_3867, SV2V_UNCONNECTED_3868, SV2V_UNCONNECTED_3869, SV2V_UNCONNECTED_3870, SV2V_UNCONNECTED_3871, SV2V_UNCONNECTED_3872, SV2V_UNCONNECTED_3873, SV2V_UNCONNECTED_3874, SV2V_UNCONNECTED_3875, SV2V_UNCONNECTED_3876, SV2V_UNCONNECTED_3877, SV2V_UNCONNECTED_3878, SV2V_UNCONNECTED_3879, SV2V_UNCONNECTED_3880, SV2V_UNCONNECTED_3881, SV2V_UNCONNECTED_3882, SV2V_UNCONNECTED_3883, SV2V_UNCONNECTED_3884, SV2V_UNCONNECTED_3885, SV2V_UNCONNECTED_3886, SV2V_UNCONNECTED_3887, SV2V_UNCONNECTED_3888, SV2V_UNCONNECTED_3889, SV2V_UNCONNECTED_3890, SV2V_UNCONNECTED_3891, SV2V_UNCONNECTED_3892, SV2V_UNCONNECTED_3893, SV2V_UNCONNECTED_3894, SV2V_UNCONNECTED_3895, SV2V_UNCONNECTED_3896, SV2V_UNCONNECTED_3897, SV2V_UNCONNECTED_3898, SV2V_UNCONNECTED_3899, SV2V_UNCONNECTED_3900, SV2V_UNCONNECTED_3901, SV2V_UNCONNECTED_3902, SV2V_UNCONNECTED_3903, SV2V_UNCONNECTED_3904, SV2V_UNCONNECTED_3905, SV2V_UNCONNECTED_3906, SV2V_UNCONNECTED_3907, SV2V_UNCONNECTED_3908, SV2V_UNCONNECTED_3909, SV2V_UNCONNECTED_3910, SV2V_UNCONNECTED_3911, SV2V_UNCONNECTED_3912, SV2V_UNCONNECTED_3913, SV2V_UNCONNECTED_3914, SV2V_UNCONNECTED_3915, SV2V_UNCONNECTED_3916, SV2V_UNCONNECTED_3917, SV2V_UNCONNECTED_3918, SV2V_UNCONNECTED_3919, SV2V_UNCONNECTED_3920, SV2V_UNCONNECTED_3921, SV2V_UNCONNECTED_3922, SV2V_UNCONNECTED_3923, SV2V_UNCONNECTED_3924, SV2V_UNCONNECTED_3925, SV2V_UNCONNECTED_3926, SV2V_UNCONNECTED_3927, SV2V_UNCONNECTED_3928, SV2V_UNCONNECTED_3929, SV2V_UNCONNECTED_3930, SV2V_UNCONNECTED_3931, SV2V_UNCONNECTED_3932, SV2V_UNCONNECTED_3933, SV2V_UNCONNECTED_3934, SV2V_UNCONNECTED_3935, SV2V_UNCONNECTED_3936, SV2V_UNCONNECTED_3937, SV2V_UNCONNECTED_3938, SV2V_UNCONNECTED_3939, SV2V_UNCONNECTED_3940, SV2V_UNCONNECTED_3941, SV2V_UNCONNECTED_3942, SV2V_UNCONNECTED_3943, SV2V_UNCONNECTED_3944, SV2V_UNCONNECTED_3945, SV2V_UNCONNECTED_3946, SV2V_UNCONNECTED_3947, SV2V_UNCONNECTED_3948, SV2V_UNCONNECTED_3949, SV2V_UNCONNECTED_3950, SV2V_UNCONNECTED_3951, SV2V_UNCONNECTED_3952, SV2V_UNCONNECTED_3953, SV2V_UNCONNECTED_3954, SV2V_UNCONNECTED_3955, SV2V_UNCONNECTED_3956, SV2V_UNCONNECTED_3957, SV2V_UNCONNECTED_3958, SV2V_UNCONNECTED_3959, SV2V_UNCONNECTED_3960, SV2V_UNCONNECTED_3961, SV2V_UNCONNECTED_3962, SV2V_UNCONNECTED_3963, SV2V_UNCONNECTED_3964, SV2V_UNCONNECTED_3965, SV2V_UNCONNECTED_3966, SV2V_UNCONNECTED_3967, SV2V_UNCONNECTED_3968, SV2V_UNCONNECTED_3969, SV2V_UNCONNECTED_3970, SV2V_UNCONNECTED_3971, SV2V_UNCONNECTED_3972, SV2V_UNCONNECTED_3973, SV2V_UNCONNECTED_3974, SV2V_UNCONNECTED_3975, SV2V_UNCONNECTED_3976, SV2V_UNCONNECTED_3977, SV2V_UNCONNECTED_3978, SV2V_UNCONNECTED_3979, SV2V_UNCONNECTED_3980, SV2V_UNCONNECTED_3981, SV2V_UNCONNECTED_3982, SV2V_UNCONNECTED_3983, SV2V_UNCONNECTED_3984, SV2V_UNCONNECTED_3985, SV2V_UNCONNECTED_3986, SV2V_UNCONNECTED_3987, SV2V_UNCONNECTED_3988, SV2V_UNCONNECTED_3989, SV2V_UNCONNECTED_3990, SV2V_UNCONNECTED_3991, SV2V_UNCONNECTED_3992, SV2V_UNCONNECTED_3993, SV2V_UNCONNECTED_3994, SV2V_UNCONNECTED_3995, SV2V_UNCONNECTED_3996, SV2V_UNCONNECTED_3997, SV2V_UNCONNECTED_3998, SV2V_UNCONNECTED_3999, SV2V_UNCONNECTED_4000, SV2V_UNCONNECTED_4001, SV2V_UNCONNECTED_4002, SV2V_UNCONNECTED_4003, SV2V_UNCONNECTED_4004, SV2V_UNCONNECTED_4005, SV2V_UNCONNECTED_4006, SV2V_UNCONNECTED_4007, SV2V_UNCONNECTED_4008, SV2V_UNCONNECTED_4009, SV2V_UNCONNECTED_4010, SV2V_UNCONNECTED_4011, SV2V_UNCONNECTED_4012, SV2V_UNCONNECTED_4013, SV2V_UNCONNECTED_4014, SV2V_UNCONNECTED_4015, SV2V_UNCONNECTED_4016, SV2V_UNCONNECTED_4017, SV2V_UNCONNECTED_4018, SV2V_UNCONNECTED_4019, SV2V_UNCONNECTED_4020, SV2V_UNCONNECTED_4021, SV2V_UNCONNECTED_4022, SV2V_UNCONNECTED_4023, SV2V_UNCONNECTED_4024, SV2V_UNCONNECTED_4025, SV2V_UNCONNECTED_4026, SV2V_UNCONNECTED_4027, SV2V_UNCONNECTED_4028, SV2V_UNCONNECTED_4029, SV2V_UNCONNECTED_4030, SV2V_UNCONNECTED_4031, SV2V_UNCONNECTED_4032, SV2V_UNCONNECTED_4033, SV2V_UNCONNECTED_4034, SV2V_UNCONNECTED_4035, SV2V_UNCONNECTED_4036, SV2V_UNCONNECTED_4037, SV2V_UNCONNECTED_4038, SV2V_UNCONNECTED_4039, SV2V_UNCONNECTED_4040, SV2V_UNCONNECTED_4041, SV2V_UNCONNECTED_4042, SV2V_UNCONNECTED_4043, SV2V_UNCONNECTED_4044, SV2V_UNCONNECTED_4045, SV2V_UNCONNECTED_4046, SV2V_UNCONNECTED_4047, SV2V_UNCONNECTED_4048, SV2V_UNCONNECTED_4049, SV2V_UNCONNECTED_4050, SV2V_UNCONNECTED_4051, SV2V_UNCONNECTED_4052, SV2V_UNCONNECTED_4053, SV2V_UNCONNECTED_4054, SV2V_UNCONNECTED_4055, SV2V_UNCONNECTED_4056, SV2V_UNCONNECTED_4057, SV2V_UNCONNECTED_4058, SV2V_UNCONNECTED_4059, SV2V_UNCONNECTED_4060, SV2V_UNCONNECTED_4061, SV2V_UNCONNECTED_4062, SV2V_UNCONNECTED_4063, SV2V_UNCONNECTED_4064, SV2V_UNCONNECTED_4065, SV2V_UNCONNECTED_4066, SV2V_UNCONNECTED_4067, SV2V_UNCONNECTED_4068, SV2V_UNCONNECTED_4069, SV2V_UNCONNECTED_4070, SV2V_UNCONNECTED_4071, SV2V_UNCONNECTED_4072, SV2V_UNCONNECTED_4073, SV2V_UNCONNECTED_4074, SV2V_UNCONNECTED_4075, SV2V_UNCONNECTED_4076, SV2V_UNCONNECTED_4077, SV2V_UNCONNECTED_4078, SV2V_UNCONNECTED_4079, SV2V_UNCONNECTED_4080, SV2V_UNCONNECTED_4081, SV2V_UNCONNECTED_4082, SV2V_UNCONNECTED_4083, SV2V_UNCONNECTED_4084, SV2V_UNCONNECTED_4085, SV2V_UNCONNECTED_4086, SV2V_UNCONNECTED_4087, SV2V_UNCONNECTED_4088, SV2V_UNCONNECTED_4089, SV2V_UNCONNECTED_4090, SV2V_UNCONNECTED_4091, SV2V_UNCONNECTED_4092, SV2V_UNCONNECTED_4093, SV2V_UNCONNECTED_4094, SV2V_UNCONNECTED_4095, SV2V_UNCONNECTED_4096, SV2V_UNCONNECTED_4097, SV2V_UNCONNECTED_4098, SV2V_UNCONNECTED_4099, SV2V_UNCONNECTED_4100, SV2V_UNCONNECTED_4101, SV2V_UNCONNECTED_4102, SV2V_UNCONNECTED_4103, SV2V_UNCONNECTED_4104, SV2V_UNCONNECTED_4105, SV2V_UNCONNECTED_4106, SV2V_UNCONNECTED_4107, SV2V_UNCONNECTED_4108, SV2V_UNCONNECTED_4109, SV2V_UNCONNECTED_4110, SV2V_UNCONNECTED_4111, SV2V_UNCONNECTED_4112, SV2V_UNCONNECTED_4113, SV2V_UNCONNECTED_4114, SV2V_UNCONNECTED_4115, SV2V_UNCONNECTED_4116, SV2V_UNCONNECTED_4117, SV2V_UNCONNECTED_4118, SV2V_UNCONNECTED_4119, SV2V_UNCONNECTED_4120, SV2V_UNCONNECTED_4121, SV2V_UNCONNECTED_4122, SV2V_UNCONNECTED_4123, SV2V_UNCONNECTED_4124, SV2V_UNCONNECTED_4125, SV2V_UNCONNECTED_4126, SV2V_UNCONNECTED_4127, SV2V_UNCONNECTED_4128, SV2V_UNCONNECTED_4129, SV2V_UNCONNECTED_4130, SV2V_UNCONNECTED_4131, SV2V_UNCONNECTED_4132, SV2V_UNCONNECTED_4133, SV2V_UNCONNECTED_4134, SV2V_UNCONNECTED_4135, SV2V_UNCONNECTED_4136, SV2V_UNCONNECTED_4137, SV2V_UNCONNECTED_4138, SV2V_UNCONNECTED_4139, SV2V_UNCONNECTED_4140, SV2V_UNCONNECTED_4141, SV2V_UNCONNECTED_4142, SV2V_UNCONNECTED_4143, SV2V_UNCONNECTED_4144, SV2V_UNCONNECTED_4145, SV2V_UNCONNECTED_4146, SV2V_UNCONNECTED_4147, SV2V_UNCONNECTED_4148, SV2V_UNCONNECTED_4149, SV2V_UNCONNECTED_4150, SV2V_UNCONNECTED_4151, SV2V_UNCONNECTED_4152, SV2V_UNCONNECTED_4153, SV2V_UNCONNECTED_4154, SV2V_UNCONNECTED_4155, SV2V_UNCONNECTED_4156, SV2V_UNCONNECTED_4157, SV2V_UNCONNECTED_4158, SV2V_UNCONNECTED_4159, SV2V_UNCONNECTED_4160, SV2V_UNCONNECTED_4161, SV2V_UNCONNECTED_4162, SV2V_UNCONNECTED_4163, SV2V_UNCONNECTED_4164, SV2V_UNCONNECTED_4165, SV2V_UNCONNECTED_4166, SV2V_UNCONNECTED_4167, SV2V_UNCONNECTED_4168, SV2V_UNCONNECTED_4169, SV2V_UNCONNECTED_4170, SV2V_UNCONNECTED_4171, SV2V_UNCONNECTED_4172, SV2V_UNCONNECTED_4173, SV2V_UNCONNECTED_4174, SV2V_UNCONNECTED_4175, SV2V_UNCONNECTED_4176, SV2V_UNCONNECTED_4177, SV2V_UNCONNECTED_4178, SV2V_UNCONNECTED_4179, SV2V_UNCONNECTED_4180, SV2V_UNCONNECTED_4181, SV2V_UNCONNECTED_4182, SV2V_UNCONNECTED_4183, SV2V_UNCONNECTED_4184, SV2V_UNCONNECTED_4185, SV2V_UNCONNECTED_4186, SV2V_UNCONNECTED_4187, SV2V_UNCONNECTED_4188, SV2V_UNCONNECTED_4189, SV2V_UNCONNECTED_4190, SV2V_UNCONNECTED_4191, SV2V_UNCONNECTED_4192, SV2V_UNCONNECTED_4193, SV2V_UNCONNECTED_4194, SV2V_UNCONNECTED_4195, SV2V_UNCONNECTED_4196, SV2V_UNCONNECTED_4197, SV2V_UNCONNECTED_4198, SV2V_UNCONNECTED_4199, SV2V_UNCONNECTED_4200, SV2V_UNCONNECTED_4201, SV2V_UNCONNECTED_4202, SV2V_UNCONNECTED_4203, SV2V_UNCONNECTED_4204, SV2V_UNCONNECTED_4205, SV2V_UNCONNECTED_4206, SV2V_UNCONNECTED_4207, SV2V_UNCONNECTED_4208, SV2V_UNCONNECTED_4209, SV2V_UNCONNECTED_4210, SV2V_UNCONNECTED_4211, SV2V_UNCONNECTED_4212, SV2V_UNCONNECTED_4213, SV2V_UNCONNECTED_4214, SV2V_UNCONNECTED_4215, SV2V_UNCONNECTED_4216, SV2V_UNCONNECTED_4217, SV2V_UNCONNECTED_4218, SV2V_UNCONNECTED_4219, SV2V_UNCONNECTED_4220, SV2V_UNCONNECTED_4221, SV2V_UNCONNECTED_4222, SV2V_UNCONNECTED_4223, SV2V_UNCONNECTED_4224, SV2V_UNCONNECTED_4225, SV2V_UNCONNECTED_4226, SV2V_UNCONNECTED_4227, SV2V_UNCONNECTED_4228, SV2V_UNCONNECTED_4229, SV2V_UNCONNECTED_4230, SV2V_UNCONNECTED_4231, SV2V_UNCONNECTED_4232, SV2V_UNCONNECTED_4233, SV2V_UNCONNECTED_4234, SV2V_UNCONNECTED_4235, SV2V_UNCONNECTED_4236, SV2V_UNCONNECTED_4237, SV2V_UNCONNECTED_4238, SV2V_UNCONNECTED_4239, SV2V_UNCONNECTED_4240, SV2V_UNCONNECTED_4241, SV2V_UNCONNECTED_4242, SV2V_UNCONNECTED_4243, SV2V_UNCONNECTED_4244, SV2V_UNCONNECTED_4245, SV2V_UNCONNECTED_4246, SV2V_UNCONNECTED_4247, SV2V_UNCONNECTED_4248, SV2V_UNCONNECTED_4249, SV2V_UNCONNECTED_4250, SV2V_UNCONNECTED_4251, SV2V_UNCONNECTED_4252, SV2V_UNCONNECTED_4253, SV2V_UNCONNECTED_4254, SV2V_UNCONNECTED_4255, SV2V_UNCONNECTED_4256, SV2V_UNCONNECTED_4257, SV2V_UNCONNECTED_4258, SV2V_UNCONNECTED_4259, SV2V_UNCONNECTED_4260, SV2V_UNCONNECTED_4261, SV2V_UNCONNECTED_4262, SV2V_UNCONNECTED_4263, SV2V_UNCONNECTED_4264, SV2V_UNCONNECTED_4265, SV2V_UNCONNECTED_4266, SV2V_UNCONNECTED_4267, SV2V_UNCONNECTED_4268, SV2V_UNCONNECTED_4269, SV2V_UNCONNECTED_4270, SV2V_UNCONNECTED_4271, SV2V_UNCONNECTED_4272, SV2V_UNCONNECTED_4273, SV2V_UNCONNECTED_4274, SV2V_UNCONNECTED_4275, SV2V_UNCONNECTED_4276, SV2V_UNCONNECTED_4277, SV2V_UNCONNECTED_4278, SV2V_UNCONNECTED_4279, SV2V_UNCONNECTED_4280, SV2V_UNCONNECTED_4281, SV2V_UNCONNECTED_4282, SV2V_UNCONNECTED_4283, SV2V_UNCONNECTED_4284, SV2V_UNCONNECTED_4285, SV2V_UNCONNECTED_4286, SV2V_UNCONNECTED_4287, SV2V_UNCONNECTED_4288, SV2V_UNCONNECTED_4289, SV2V_UNCONNECTED_4290, SV2V_UNCONNECTED_4291, SV2V_UNCONNECTED_4292, SV2V_UNCONNECTED_4293, SV2V_UNCONNECTED_4294, SV2V_UNCONNECTED_4295, SV2V_UNCONNECTED_4296, SV2V_UNCONNECTED_4297, SV2V_UNCONNECTED_4298, SV2V_UNCONNECTED_4299, SV2V_UNCONNECTED_4300, SV2V_UNCONNECTED_4301, SV2V_UNCONNECTED_4302, SV2V_UNCONNECTED_4303, SV2V_UNCONNECTED_4304, SV2V_UNCONNECTED_4305, SV2V_UNCONNECTED_4306, SV2V_UNCONNECTED_4307, SV2V_UNCONNECTED_4308, SV2V_UNCONNECTED_4309, SV2V_UNCONNECTED_4310, SV2V_UNCONNECTED_4311, SV2V_UNCONNECTED_4312, SV2V_UNCONNECTED_4313, SV2V_UNCONNECTED_4314, SV2V_UNCONNECTED_4315, SV2V_UNCONNECTED_4316, SV2V_UNCONNECTED_4317, SV2V_UNCONNECTED_4318, SV2V_UNCONNECTED_4319, SV2V_UNCONNECTED_4320, SV2V_UNCONNECTED_4321, SV2V_UNCONNECTED_4322, SV2V_UNCONNECTED_4323, SV2V_UNCONNECTED_4324, SV2V_UNCONNECTED_4325, SV2V_UNCONNECTED_4326, SV2V_UNCONNECTED_4327, SV2V_UNCONNECTED_4328, SV2V_UNCONNECTED_4329, SV2V_UNCONNECTED_4330, SV2V_UNCONNECTED_4331, SV2V_UNCONNECTED_4332, SV2V_UNCONNECTED_4333, SV2V_UNCONNECTED_4334, SV2V_UNCONNECTED_4335, SV2V_UNCONNECTED_4336, SV2V_UNCONNECTED_4337, SV2V_UNCONNECTED_4338, SV2V_UNCONNECTED_4339, SV2V_UNCONNECTED_4340, SV2V_UNCONNECTED_4341, SV2V_UNCONNECTED_4342, SV2V_UNCONNECTED_4343, SV2V_UNCONNECTED_4344, SV2V_UNCONNECTED_4345, SV2V_UNCONNECTED_4346, SV2V_UNCONNECTED_4347, SV2V_UNCONNECTED_4348, SV2V_UNCONNECTED_4349, SV2V_UNCONNECTED_4350, SV2V_UNCONNECTED_4351, SV2V_UNCONNECTED_4352, SV2V_UNCONNECTED_4353, SV2V_UNCONNECTED_4354, SV2V_UNCONNECTED_4355, SV2V_UNCONNECTED_4356, SV2V_UNCONNECTED_4357, SV2V_UNCONNECTED_4358, SV2V_UNCONNECTED_4359, SV2V_UNCONNECTED_4360, SV2V_UNCONNECTED_4361, SV2V_UNCONNECTED_4362, SV2V_UNCONNECTED_4363, SV2V_UNCONNECTED_4364, SV2V_UNCONNECTED_4365, SV2V_UNCONNECTED_4366, SV2V_UNCONNECTED_4367, SV2V_UNCONNECTED_4368, SV2V_UNCONNECTED_4369, SV2V_UNCONNECTED_4370, SV2V_UNCONNECTED_4371, SV2V_UNCONNECTED_4372, SV2V_UNCONNECTED_4373, SV2V_UNCONNECTED_4374, SV2V_UNCONNECTED_4375, SV2V_UNCONNECTED_4376, SV2V_UNCONNECTED_4377, SV2V_UNCONNECTED_4378, SV2V_UNCONNECTED_4379, SV2V_UNCONNECTED_4380, SV2V_UNCONNECTED_4381, SV2V_UNCONNECTED_4382, SV2V_UNCONNECTED_4383, SV2V_UNCONNECTED_4384, SV2V_UNCONNECTED_4385, SV2V_UNCONNECTED_4386, SV2V_UNCONNECTED_4387, SV2V_UNCONNECTED_4388, SV2V_UNCONNECTED_4389, SV2V_UNCONNECTED_4390, SV2V_UNCONNECTED_4391, SV2V_UNCONNECTED_4392, SV2V_UNCONNECTED_4393, SV2V_UNCONNECTED_4394, SV2V_UNCONNECTED_4395, SV2V_UNCONNECTED_4396, SV2V_UNCONNECTED_4397, SV2V_UNCONNECTED_4398, SV2V_UNCONNECTED_4399, SV2V_UNCONNECTED_4400, SV2V_UNCONNECTED_4401, SV2V_UNCONNECTED_4402, SV2V_UNCONNECTED_4403, SV2V_UNCONNECTED_4404, SV2V_UNCONNECTED_4405, SV2V_UNCONNECTED_4406, SV2V_UNCONNECTED_4407, SV2V_UNCONNECTED_4408, SV2V_UNCONNECTED_4409, SV2V_UNCONNECTED_4410, SV2V_UNCONNECTED_4411, SV2V_UNCONNECTED_4412, SV2V_UNCONNECTED_4413, SV2V_UNCONNECTED_4414, SV2V_UNCONNECTED_4415, SV2V_UNCONNECTED_4416, SV2V_UNCONNECTED_4417, SV2V_UNCONNECTED_4418, SV2V_UNCONNECTED_4419, SV2V_UNCONNECTED_4420, SV2V_UNCONNECTED_4421, SV2V_UNCONNECTED_4422, SV2V_UNCONNECTED_4423, SV2V_UNCONNECTED_4424, SV2V_UNCONNECTED_4425, SV2V_UNCONNECTED_4426, SV2V_UNCONNECTED_4427, SV2V_UNCONNECTED_4428, SV2V_UNCONNECTED_4429, SV2V_UNCONNECTED_4430, SV2V_UNCONNECTED_4431, SV2V_UNCONNECTED_4432, SV2V_UNCONNECTED_4433, SV2V_UNCONNECTED_4434, SV2V_UNCONNECTED_4435, SV2V_UNCONNECTED_4436, SV2V_UNCONNECTED_4437, SV2V_UNCONNECTED_4438, SV2V_UNCONNECTED_4439, SV2V_UNCONNECTED_4440, SV2V_UNCONNECTED_4441, SV2V_UNCONNECTED_4442, SV2V_UNCONNECTED_4443, SV2V_UNCONNECTED_4444, SV2V_UNCONNECTED_4445, SV2V_UNCONNECTED_4446, SV2V_UNCONNECTED_4447, SV2V_UNCONNECTED_4448, SV2V_UNCONNECTED_4449, SV2V_UNCONNECTED_4450, SV2V_UNCONNECTED_4451, SV2V_UNCONNECTED_4452, SV2V_UNCONNECTED_4453, SV2V_UNCONNECTED_4454, SV2V_UNCONNECTED_4455, SV2V_UNCONNECTED_4456, SV2V_UNCONNECTED_4457, SV2V_UNCONNECTED_4458, SV2V_UNCONNECTED_4459, SV2V_UNCONNECTED_4460, SV2V_UNCONNECTED_4461, SV2V_UNCONNECTED_4462, SV2V_UNCONNECTED_4463, SV2V_UNCONNECTED_4464, SV2V_UNCONNECTED_4465, SV2V_UNCONNECTED_4466, SV2V_UNCONNECTED_4467, SV2V_UNCONNECTED_4468, SV2V_UNCONNECTED_4469, SV2V_UNCONNECTED_4470, SV2V_UNCONNECTED_4471, SV2V_UNCONNECTED_4472, SV2V_UNCONNECTED_4473, SV2V_UNCONNECTED_4474, SV2V_UNCONNECTED_4475, SV2V_UNCONNECTED_4476, SV2V_UNCONNECTED_4477, SV2V_UNCONNECTED_4478, SV2V_UNCONNECTED_4479, SV2V_UNCONNECTED_4480, SV2V_UNCONNECTED_4481, SV2V_UNCONNECTED_4482, SV2V_UNCONNECTED_4483, SV2V_UNCONNECTED_4484, SV2V_UNCONNECTED_4485, SV2V_UNCONNECTED_4486, SV2V_UNCONNECTED_4487, SV2V_UNCONNECTED_4488, SV2V_UNCONNECTED_4489, SV2V_UNCONNECTED_4490, SV2V_UNCONNECTED_4491, SV2V_UNCONNECTED_4492, SV2V_UNCONNECTED_4493, SV2V_UNCONNECTED_4494, SV2V_UNCONNECTED_4495, SV2V_UNCONNECTED_4496, SV2V_UNCONNECTED_4497, SV2V_UNCONNECTED_4498, SV2V_UNCONNECTED_4499, SV2V_UNCONNECTED_4500, SV2V_UNCONNECTED_4501, SV2V_UNCONNECTED_4502, SV2V_UNCONNECTED_4503, SV2V_UNCONNECTED_4504, SV2V_UNCONNECTED_4505, SV2V_UNCONNECTED_4506, SV2V_UNCONNECTED_4507, SV2V_UNCONNECTED_4508, SV2V_UNCONNECTED_4509, SV2V_UNCONNECTED_4510, SV2V_UNCONNECTED_4511, SV2V_UNCONNECTED_4512, SV2V_UNCONNECTED_4513, SV2V_UNCONNECTED_4514, SV2V_UNCONNECTED_4515, SV2V_UNCONNECTED_4516, SV2V_UNCONNECTED_4517, SV2V_UNCONNECTED_4518, SV2V_UNCONNECTED_4519, SV2V_UNCONNECTED_4520, SV2V_UNCONNECTED_4521, SV2V_UNCONNECTED_4522, SV2V_UNCONNECTED_4523, SV2V_UNCONNECTED_4524, SV2V_UNCONNECTED_4525, SV2V_UNCONNECTED_4526, SV2V_UNCONNECTED_4527, SV2V_UNCONNECTED_4528, SV2V_UNCONNECTED_4529, SV2V_UNCONNECTED_4530, SV2V_UNCONNECTED_4531, SV2V_UNCONNECTED_4532, SV2V_UNCONNECTED_4533, SV2V_UNCONNECTED_4534, SV2V_UNCONNECTED_4535, SV2V_UNCONNECTED_4536, SV2V_UNCONNECTED_4537, SV2V_UNCONNECTED_4538, SV2V_UNCONNECTED_4539, SV2V_UNCONNECTED_4540, SV2V_UNCONNECTED_4541, SV2V_UNCONNECTED_4542, SV2V_UNCONNECTED_4543, SV2V_UNCONNECTED_4544, SV2V_UNCONNECTED_4545, SV2V_UNCONNECTED_4546, SV2V_UNCONNECTED_4547, SV2V_UNCONNECTED_4548, SV2V_UNCONNECTED_4549, SV2V_UNCONNECTED_4550, SV2V_UNCONNECTED_4551, SV2V_UNCONNECTED_4552, SV2V_UNCONNECTED_4553, SV2V_UNCONNECTED_4554, SV2V_UNCONNECTED_4555, SV2V_UNCONNECTED_4556, SV2V_UNCONNECTED_4557, SV2V_UNCONNECTED_4558, SV2V_UNCONNECTED_4559, SV2V_UNCONNECTED_4560, SV2V_UNCONNECTED_4561, SV2V_UNCONNECTED_4562, SV2V_UNCONNECTED_4563, SV2V_UNCONNECTED_4564, SV2V_UNCONNECTED_4565, SV2V_UNCONNECTED_4566, SV2V_UNCONNECTED_4567, SV2V_UNCONNECTED_4568, SV2V_UNCONNECTED_4569, SV2V_UNCONNECTED_4570, SV2V_UNCONNECTED_4571, SV2V_UNCONNECTED_4572, SV2V_UNCONNECTED_4573, SV2V_UNCONNECTED_4574, SV2V_UNCONNECTED_4575, SV2V_UNCONNECTED_4576, SV2V_UNCONNECTED_4577, SV2V_UNCONNECTED_4578, SV2V_UNCONNECTED_4579, SV2V_UNCONNECTED_4580, SV2V_UNCONNECTED_4581, SV2V_UNCONNECTED_4582, SV2V_UNCONNECTED_4583, SV2V_UNCONNECTED_4584, SV2V_UNCONNECTED_4585, SV2V_UNCONNECTED_4586, SV2V_UNCONNECTED_4587, SV2V_UNCONNECTED_4588, SV2V_UNCONNECTED_4589, SV2V_UNCONNECTED_4590, SV2V_UNCONNECTED_4591, SV2V_UNCONNECTED_4592, SV2V_UNCONNECTED_4593, SV2V_UNCONNECTED_4594, SV2V_UNCONNECTED_4595, SV2V_UNCONNECTED_4596, SV2V_UNCONNECTED_4597, SV2V_UNCONNECTED_4598, SV2V_UNCONNECTED_4599, SV2V_UNCONNECTED_4600, SV2V_UNCONNECTED_4601, SV2V_UNCONNECTED_4602, SV2V_UNCONNECTED_4603, SV2V_UNCONNECTED_4604, SV2V_UNCONNECTED_4605, SV2V_UNCONNECTED_4606, SV2V_UNCONNECTED_4607, SV2V_UNCONNECTED_4608, SV2V_UNCONNECTED_4609, SV2V_UNCONNECTED_4610, SV2V_UNCONNECTED_4611, SV2V_UNCONNECTED_4612, SV2V_UNCONNECTED_4613, SV2V_UNCONNECTED_4614, SV2V_UNCONNECTED_4615, SV2V_UNCONNECTED_4616, SV2V_UNCONNECTED_4617, SV2V_UNCONNECTED_4618, SV2V_UNCONNECTED_4619, SV2V_UNCONNECTED_4620, SV2V_UNCONNECTED_4621, SV2V_UNCONNECTED_4622, SV2V_UNCONNECTED_4623, SV2V_UNCONNECTED_4624, SV2V_UNCONNECTED_4625, SV2V_UNCONNECTED_4626, SV2V_UNCONNECTED_4627, SV2V_UNCONNECTED_4628, SV2V_UNCONNECTED_4629, SV2V_UNCONNECTED_4630, SV2V_UNCONNECTED_4631, SV2V_UNCONNECTED_4632, SV2V_UNCONNECTED_4633, SV2V_UNCONNECTED_4634, SV2V_UNCONNECTED_4635, SV2V_UNCONNECTED_4636, SV2V_UNCONNECTED_4637, SV2V_UNCONNECTED_4638, SV2V_UNCONNECTED_4639, SV2V_UNCONNECTED_4640, SV2V_UNCONNECTED_4641, SV2V_UNCONNECTED_4642, SV2V_UNCONNECTED_4643, SV2V_UNCONNECTED_4644, SV2V_UNCONNECTED_4645, SV2V_UNCONNECTED_4646, SV2V_UNCONNECTED_4647, SV2V_UNCONNECTED_4648, SV2V_UNCONNECTED_4649, SV2V_UNCONNECTED_4650, SV2V_UNCONNECTED_4651, SV2V_UNCONNECTED_4652, SV2V_UNCONNECTED_4653, SV2V_UNCONNECTED_4654, SV2V_UNCONNECTED_4655, SV2V_UNCONNECTED_4656, SV2V_UNCONNECTED_4657, SV2V_UNCONNECTED_4658, SV2V_UNCONNECTED_4659, SV2V_UNCONNECTED_4660, SV2V_UNCONNECTED_4661, SV2V_UNCONNECTED_4662, SV2V_UNCONNECTED_4663, SV2V_UNCONNECTED_4664, SV2V_UNCONNECTED_4665, SV2V_UNCONNECTED_4666, SV2V_UNCONNECTED_4667, SV2V_UNCONNECTED_4668, SV2V_UNCONNECTED_4669, SV2V_UNCONNECTED_4670, SV2V_UNCONNECTED_4671, SV2V_UNCONNECTED_4672, SV2V_UNCONNECTED_4673, SV2V_UNCONNECTED_4674, SV2V_UNCONNECTED_4675, SV2V_UNCONNECTED_4676, SV2V_UNCONNECTED_4677, SV2V_UNCONNECTED_4678, SV2V_UNCONNECTED_4679, SV2V_UNCONNECTED_4680, SV2V_UNCONNECTED_4681, SV2V_UNCONNECTED_4682, SV2V_UNCONNECTED_4683, SV2V_UNCONNECTED_4684, SV2V_UNCONNECTED_4685, SV2V_UNCONNECTED_4686, SV2V_UNCONNECTED_4687, SV2V_UNCONNECTED_4688, SV2V_UNCONNECTED_4689, SV2V_UNCONNECTED_4690, SV2V_UNCONNECTED_4691, SV2V_UNCONNECTED_4692, SV2V_UNCONNECTED_4693, SV2V_UNCONNECTED_4694, SV2V_UNCONNECTED_4695, SV2V_UNCONNECTED_4696, SV2V_UNCONNECTED_4697, SV2V_UNCONNECTED_4698, SV2V_UNCONNECTED_4699, SV2V_UNCONNECTED_4700, SV2V_UNCONNECTED_4701, SV2V_UNCONNECTED_4702, SV2V_UNCONNECTED_4703, SV2V_UNCONNECTED_4704, SV2V_UNCONNECTED_4705, SV2V_UNCONNECTED_4706, SV2V_UNCONNECTED_4707, SV2V_UNCONNECTED_4708, SV2V_UNCONNECTED_4709, SV2V_UNCONNECTED_4710, SV2V_UNCONNECTED_4711, SV2V_UNCONNECTED_4712, SV2V_UNCONNECTED_4713, SV2V_UNCONNECTED_4714, SV2V_UNCONNECTED_4715, SV2V_UNCONNECTED_4716, SV2V_UNCONNECTED_4717, SV2V_UNCONNECTED_4718, SV2V_UNCONNECTED_4719, SV2V_UNCONNECTED_4720, SV2V_UNCONNECTED_4721, SV2V_UNCONNECTED_4722, SV2V_UNCONNECTED_4723, SV2V_UNCONNECTED_4724, SV2V_UNCONNECTED_4725, SV2V_UNCONNECTED_4726, SV2V_UNCONNECTED_4727, SV2V_UNCONNECTED_4728, SV2V_UNCONNECTED_4729, SV2V_UNCONNECTED_4730, SV2V_UNCONNECTED_4731, SV2V_UNCONNECTED_4732, SV2V_UNCONNECTED_4733, SV2V_UNCONNECTED_4734, SV2V_UNCONNECTED_4735, SV2V_UNCONNECTED_4736, SV2V_UNCONNECTED_4737, SV2V_UNCONNECTED_4738, SV2V_UNCONNECTED_4739, SV2V_UNCONNECTED_4740, SV2V_UNCONNECTED_4741, SV2V_UNCONNECTED_4742, SV2V_UNCONNECTED_4743, SV2V_UNCONNECTED_4744, SV2V_UNCONNECTED_4745, SV2V_UNCONNECTED_4746, SV2V_UNCONNECTED_4747, SV2V_UNCONNECTED_4748, SV2V_UNCONNECTED_4749, SV2V_UNCONNECTED_4750, SV2V_UNCONNECTED_4751, SV2V_UNCONNECTED_4752, SV2V_UNCONNECTED_4753, SV2V_UNCONNECTED_4754, SV2V_UNCONNECTED_4755, SV2V_UNCONNECTED_4756, SV2V_UNCONNECTED_4757, SV2V_UNCONNECTED_4758, SV2V_UNCONNECTED_4759, SV2V_UNCONNECTED_4760, SV2V_UNCONNECTED_4761, SV2V_UNCONNECTED_4762, SV2V_UNCONNECTED_4763, SV2V_UNCONNECTED_4764, SV2V_UNCONNECTED_4765, SV2V_UNCONNECTED_4766, SV2V_UNCONNECTED_4767, SV2V_UNCONNECTED_4768, SV2V_UNCONNECTED_4769, SV2V_UNCONNECTED_4770, SV2V_UNCONNECTED_4771, SV2V_UNCONNECTED_4772, SV2V_UNCONNECTED_4773, SV2V_UNCONNECTED_4774, SV2V_UNCONNECTED_4775, SV2V_UNCONNECTED_4776, SV2V_UNCONNECTED_4777, SV2V_UNCONNECTED_4778, SV2V_UNCONNECTED_4779, SV2V_UNCONNECTED_4780, SV2V_UNCONNECTED_4781, SV2V_UNCONNECTED_4782, SV2V_UNCONNECTED_4783, SV2V_UNCONNECTED_4784, SV2V_UNCONNECTED_4785, SV2V_UNCONNECTED_4786, SV2V_UNCONNECTED_4787, SV2V_UNCONNECTED_4788, SV2V_UNCONNECTED_4789, SV2V_UNCONNECTED_4790, SV2V_UNCONNECTED_4791, SV2V_UNCONNECTED_4792, SV2V_UNCONNECTED_4793, SV2V_UNCONNECTED_4794, SV2V_UNCONNECTED_4795, SV2V_UNCONNECTED_4796, SV2V_UNCONNECTED_4797, SV2V_UNCONNECTED_4798, SV2V_UNCONNECTED_4799, SV2V_UNCONNECTED_4800, SV2V_UNCONNECTED_4801, SV2V_UNCONNECTED_4802, SV2V_UNCONNECTED_4803, SV2V_UNCONNECTED_4804, SV2V_UNCONNECTED_4805, SV2V_UNCONNECTED_4806, SV2V_UNCONNECTED_4807, SV2V_UNCONNECTED_4808, SV2V_UNCONNECTED_4809, SV2V_UNCONNECTED_4810, SV2V_UNCONNECTED_4811, SV2V_UNCONNECTED_4812, SV2V_UNCONNECTED_4813, SV2V_UNCONNECTED_4814, SV2V_UNCONNECTED_4815, SV2V_UNCONNECTED_4816, SV2V_UNCONNECTED_4817, SV2V_UNCONNECTED_4818, SV2V_UNCONNECTED_4819, SV2V_UNCONNECTED_4820, SV2V_UNCONNECTED_4821, SV2V_UNCONNECTED_4822, SV2V_UNCONNECTED_4823, SV2V_UNCONNECTED_4824, SV2V_UNCONNECTED_4825, SV2V_UNCONNECTED_4826, SV2V_UNCONNECTED_4827, SV2V_UNCONNECTED_4828, SV2V_UNCONNECTED_4829, SV2V_UNCONNECTED_4830, SV2V_UNCONNECTED_4831, SV2V_UNCONNECTED_4832, SV2V_UNCONNECTED_4833, SV2V_UNCONNECTED_4834, SV2V_UNCONNECTED_4835, SV2V_UNCONNECTED_4836, SV2V_UNCONNECTED_4837, SV2V_UNCONNECTED_4838, SV2V_UNCONNECTED_4839, SV2V_UNCONNECTED_4840, SV2V_UNCONNECTED_4841, SV2V_UNCONNECTED_4842, SV2V_UNCONNECTED_4843, SV2V_UNCONNECTED_4844, SV2V_UNCONNECTED_4845, SV2V_UNCONNECTED_4846, SV2V_UNCONNECTED_4847, SV2V_UNCONNECTED_4848, SV2V_UNCONNECTED_4849, SV2V_UNCONNECTED_4850, SV2V_UNCONNECTED_4851, SV2V_UNCONNECTED_4852, SV2V_UNCONNECTED_4853, SV2V_UNCONNECTED_4854, SV2V_UNCONNECTED_4855, SV2V_UNCONNECTED_4856, SV2V_UNCONNECTED_4857, SV2V_UNCONNECTED_4858, SV2V_UNCONNECTED_4859, SV2V_UNCONNECTED_4860, SV2V_UNCONNECTED_4861, SV2V_UNCONNECTED_4862, SV2V_UNCONNECTED_4863, SV2V_UNCONNECTED_4864, SV2V_UNCONNECTED_4865, SV2V_UNCONNECTED_4866, SV2V_UNCONNECTED_4867, SV2V_UNCONNECTED_4868, SV2V_UNCONNECTED_4869, SV2V_UNCONNECTED_4870, SV2V_UNCONNECTED_4871, SV2V_UNCONNECTED_4872, SV2V_UNCONNECTED_4873, SV2V_UNCONNECTED_4874, SV2V_UNCONNECTED_4875, SV2V_UNCONNECTED_4876, SV2V_UNCONNECTED_4877, SV2V_UNCONNECTED_4878, SV2V_UNCONNECTED_4879, SV2V_UNCONNECTED_4880, SV2V_UNCONNECTED_4881, SV2V_UNCONNECTED_4882, SV2V_UNCONNECTED_4883, SV2V_UNCONNECTED_4884, SV2V_UNCONNECTED_4885, SV2V_UNCONNECTED_4886, SV2V_UNCONNECTED_4887, SV2V_UNCONNECTED_4888, SV2V_UNCONNECTED_4889, SV2V_UNCONNECTED_4890, SV2V_UNCONNECTED_4891, SV2V_UNCONNECTED_4892, SV2V_UNCONNECTED_4893, SV2V_UNCONNECTED_4894, SV2V_UNCONNECTED_4895, SV2V_UNCONNECTED_4896, SV2V_UNCONNECTED_4897, SV2V_UNCONNECTED_4898, SV2V_UNCONNECTED_4899, SV2V_UNCONNECTED_4900, SV2V_UNCONNECTED_4901, SV2V_UNCONNECTED_4902, SV2V_UNCONNECTED_4903, SV2V_UNCONNECTED_4904, SV2V_UNCONNECTED_4905, SV2V_UNCONNECTED_4906, SV2V_UNCONNECTED_4907, SV2V_UNCONNECTED_4908, SV2V_UNCONNECTED_4909, SV2V_UNCONNECTED_4910, SV2V_UNCONNECTED_4911, SV2V_UNCONNECTED_4912, SV2V_UNCONNECTED_4913, SV2V_UNCONNECTED_4914, SV2V_UNCONNECTED_4915, SV2V_UNCONNECTED_4916, SV2V_UNCONNECTED_4917, SV2V_UNCONNECTED_4918, SV2V_UNCONNECTED_4919, SV2V_UNCONNECTED_4920, SV2V_UNCONNECTED_4921, SV2V_UNCONNECTED_4922, SV2V_UNCONNECTED_4923, SV2V_UNCONNECTED_4924, SV2V_UNCONNECTED_4925, SV2V_UNCONNECTED_4926, SV2V_UNCONNECTED_4927, SV2V_UNCONNECTED_4928, SV2V_UNCONNECTED_4929, SV2V_UNCONNECTED_4930, SV2V_UNCONNECTED_4931, SV2V_UNCONNECTED_4932, SV2V_UNCONNECTED_4933, SV2V_UNCONNECTED_4934, SV2V_UNCONNECTED_4935, SV2V_UNCONNECTED_4936, SV2V_UNCONNECTED_4937, SV2V_UNCONNECTED_4938, SV2V_UNCONNECTED_4939, SV2V_UNCONNECTED_4940, SV2V_UNCONNECTED_4941, SV2V_UNCONNECTED_4942, SV2V_UNCONNECTED_4943, SV2V_UNCONNECTED_4944, SV2V_UNCONNECTED_4945, SV2V_UNCONNECTED_4946, SV2V_UNCONNECTED_4947, SV2V_UNCONNECTED_4948, SV2V_UNCONNECTED_4949, SV2V_UNCONNECTED_4950, SV2V_UNCONNECTED_4951, SV2V_UNCONNECTED_4952, SV2V_UNCONNECTED_4953, SV2V_UNCONNECTED_4954, SV2V_UNCONNECTED_4955, SV2V_UNCONNECTED_4956, SV2V_UNCONNECTED_4957, SV2V_UNCONNECTED_4958, SV2V_UNCONNECTED_4959, SV2V_UNCONNECTED_4960, SV2V_UNCONNECTED_4961, SV2V_UNCONNECTED_4962, SV2V_UNCONNECTED_4963, SV2V_UNCONNECTED_4964, SV2V_UNCONNECTED_4965, SV2V_UNCONNECTED_4966, SV2V_UNCONNECTED_4967, SV2V_UNCONNECTED_4968, SV2V_UNCONNECTED_4969, SV2V_UNCONNECTED_4970, SV2V_UNCONNECTED_4971, SV2V_UNCONNECTED_4972, SV2V_UNCONNECTED_4973, SV2V_UNCONNECTED_4974, SV2V_UNCONNECTED_4975, SV2V_UNCONNECTED_4976, SV2V_UNCONNECTED_4977, SV2V_UNCONNECTED_4978, SV2V_UNCONNECTED_4979, SV2V_UNCONNECTED_4980, SV2V_UNCONNECTED_4981, SV2V_UNCONNECTED_4982, SV2V_UNCONNECTED_4983, SV2V_UNCONNECTED_4984, SV2V_UNCONNECTED_4985, SV2V_UNCONNECTED_4986, SV2V_UNCONNECTED_4987, SV2V_UNCONNECTED_4988, SV2V_UNCONNECTED_4989, SV2V_UNCONNECTED_4990, SV2V_UNCONNECTED_4991, SV2V_UNCONNECTED_4992, SV2V_UNCONNECTED_4993, SV2V_UNCONNECTED_4994, SV2V_UNCONNECTED_4995, SV2V_UNCONNECTED_4996, SV2V_UNCONNECTED_4997, SV2V_UNCONNECTED_4998, SV2V_UNCONNECTED_4999, SV2V_UNCONNECTED_5000, SV2V_UNCONNECTED_5001, SV2V_UNCONNECTED_5002, SV2V_UNCONNECTED_5003, SV2V_UNCONNECTED_5004, SV2V_UNCONNECTED_5005, SV2V_UNCONNECTED_5006, SV2V_UNCONNECTED_5007, SV2V_UNCONNECTED_5008, SV2V_UNCONNECTED_5009, SV2V_UNCONNECTED_5010, SV2V_UNCONNECTED_5011, SV2V_UNCONNECTED_5012, SV2V_UNCONNECTED_5013, SV2V_UNCONNECTED_5014, SV2V_UNCONNECTED_5015, SV2V_UNCONNECTED_5016, SV2V_UNCONNECTED_5017, SV2V_UNCONNECTED_5018, SV2V_UNCONNECTED_5019, SV2V_UNCONNECTED_5020, SV2V_UNCONNECTED_5021, SV2V_UNCONNECTED_5022, SV2V_UNCONNECTED_5023, SV2V_UNCONNECTED_5024, SV2V_UNCONNECTED_5025, SV2V_UNCONNECTED_5026, SV2V_UNCONNECTED_5027, SV2V_UNCONNECTED_5028, SV2V_UNCONNECTED_5029, SV2V_UNCONNECTED_5030, SV2V_UNCONNECTED_5031, SV2V_UNCONNECTED_5032, SV2V_UNCONNECTED_5033, SV2V_UNCONNECTED_5034, SV2V_UNCONNECTED_5035, SV2V_UNCONNECTED_5036, SV2V_UNCONNECTED_5037, SV2V_UNCONNECTED_5038, SV2V_UNCONNECTED_5039, SV2V_UNCONNECTED_5040, SV2V_UNCONNECTED_5041, SV2V_UNCONNECTED_5042, SV2V_UNCONNECTED_5043, SV2V_UNCONNECTED_5044, SV2V_UNCONNECTED_5045, SV2V_UNCONNECTED_5046, SV2V_UNCONNECTED_5047, SV2V_UNCONNECTED_5048, SV2V_UNCONNECTED_5049, SV2V_UNCONNECTED_5050, SV2V_UNCONNECTED_5051, SV2V_UNCONNECTED_5052, SV2V_UNCONNECTED_5053, SV2V_UNCONNECTED_5054, SV2V_UNCONNECTED_5055, SV2V_UNCONNECTED_5056, SV2V_UNCONNECTED_5057, SV2V_UNCONNECTED_5058, SV2V_UNCONNECTED_5059, SV2V_UNCONNECTED_5060, SV2V_UNCONNECTED_5061, SV2V_UNCONNECTED_5062, SV2V_UNCONNECTED_5063, SV2V_UNCONNECTED_5064, SV2V_UNCONNECTED_5065, SV2V_UNCONNECTED_5066, SV2V_UNCONNECTED_5067, SV2V_UNCONNECTED_5068, SV2V_UNCONNECTED_5069, SV2V_UNCONNECTED_5070, SV2V_UNCONNECTED_5071, SV2V_UNCONNECTED_5072, SV2V_UNCONNECTED_5073, SV2V_UNCONNECTED_5074, SV2V_UNCONNECTED_5075, SV2V_UNCONNECTED_5076, SV2V_UNCONNECTED_5077, SV2V_UNCONNECTED_5078, SV2V_UNCONNECTED_5079, SV2V_UNCONNECTED_5080, SV2V_UNCONNECTED_5081, SV2V_UNCONNECTED_5082, SV2V_UNCONNECTED_5083, SV2V_UNCONNECTED_5084, SV2V_UNCONNECTED_5085, SV2V_UNCONNECTED_5086, SV2V_UNCONNECTED_5087, SV2V_UNCONNECTED_5088, SV2V_UNCONNECTED_5089, SV2V_UNCONNECTED_5090, SV2V_UNCONNECTED_5091, SV2V_UNCONNECTED_5092, SV2V_UNCONNECTED_5093, SV2V_UNCONNECTED_5094, SV2V_UNCONNECTED_5095, SV2V_UNCONNECTED_5096, SV2V_UNCONNECTED_5097, SV2V_UNCONNECTED_5098, SV2V_UNCONNECTED_5099, SV2V_UNCONNECTED_5100, SV2V_UNCONNECTED_5101, SV2V_UNCONNECTED_5102, SV2V_UNCONNECTED_5103, SV2V_UNCONNECTED_5104, SV2V_UNCONNECTED_5105, SV2V_UNCONNECTED_5106, SV2V_UNCONNECTED_5107, SV2V_UNCONNECTED_5108, SV2V_UNCONNECTED_5109, SV2V_UNCONNECTED_5110, SV2V_UNCONNECTED_5111, SV2V_UNCONNECTED_5112, SV2V_UNCONNECTED_5113, SV2V_UNCONNECTED_5114, SV2V_UNCONNECTED_5115, SV2V_UNCONNECTED_5116, SV2V_UNCONNECTED_5117, SV2V_UNCONNECTED_5118, SV2V_UNCONNECTED_5119, SV2V_UNCONNECTED_5120, SV2V_UNCONNECTED_5121, SV2V_UNCONNECTED_5122, SV2V_UNCONNECTED_5123, SV2V_UNCONNECTED_5124, SV2V_UNCONNECTED_5125, SV2V_UNCONNECTED_5126, SV2V_UNCONNECTED_5127, SV2V_UNCONNECTED_5128, SV2V_UNCONNECTED_5129, SV2V_UNCONNECTED_5130, SV2V_UNCONNECTED_5131, SV2V_UNCONNECTED_5132, SV2V_UNCONNECTED_5133, SV2V_UNCONNECTED_5134, SV2V_UNCONNECTED_5135, SV2V_UNCONNECTED_5136, SV2V_UNCONNECTED_5137, SV2V_UNCONNECTED_5138, SV2V_UNCONNECTED_5139, SV2V_UNCONNECTED_5140, SV2V_UNCONNECTED_5141, SV2V_UNCONNECTED_5142, SV2V_UNCONNECTED_5143, SV2V_UNCONNECTED_5144, SV2V_UNCONNECTED_5145, SV2V_UNCONNECTED_5146, SV2V_UNCONNECTED_5147, SV2V_UNCONNECTED_5148, SV2V_UNCONNECTED_5149, SV2V_UNCONNECTED_5150, SV2V_UNCONNECTED_5151, SV2V_UNCONNECTED_5152, SV2V_UNCONNECTED_5153, SV2V_UNCONNECTED_5154, SV2V_UNCONNECTED_5155, SV2V_UNCONNECTED_5156, SV2V_UNCONNECTED_5157, SV2V_UNCONNECTED_5158, SV2V_UNCONNECTED_5159, SV2V_UNCONNECTED_5160, SV2V_UNCONNECTED_5161, SV2V_UNCONNECTED_5162, SV2V_UNCONNECTED_5163, SV2V_UNCONNECTED_5164, SV2V_UNCONNECTED_5165, SV2V_UNCONNECTED_5166, SV2V_UNCONNECTED_5167, SV2V_UNCONNECTED_5168, SV2V_UNCONNECTED_5169, SV2V_UNCONNECTED_5170, SV2V_UNCONNECTED_5171, SV2V_UNCONNECTED_5172, SV2V_UNCONNECTED_5173, SV2V_UNCONNECTED_5174, SV2V_UNCONNECTED_5175, SV2V_UNCONNECTED_5176, SV2V_UNCONNECTED_5177, SV2V_UNCONNECTED_5178, SV2V_UNCONNECTED_5179, SV2V_UNCONNECTED_5180, SV2V_UNCONNECTED_5181, SV2V_UNCONNECTED_5182, SV2V_UNCONNECTED_5183, SV2V_UNCONNECTED_5184, SV2V_UNCONNECTED_5185, SV2V_UNCONNECTED_5186, SV2V_UNCONNECTED_5187, SV2V_UNCONNECTED_5188, SV2V_UNCONNECTED_5189, SV2V_UNCONNECTED_5190, SV2V_UNCONNECTED_5191, SV2V_UNCONNECTED_5192, SV2V_UNCONNECTED_5193, SV2V_UNCONNECTED_5194, SV2V_UNCONNECTED_5195, SV2V_UNCONNECTED_5196, SV2V_UNCONNECTED_5197, SV2V_UNCONNECTED_5198, SV2V_UNCONNECTED_5199, SV2V_UNCONNECTED_5200, SV2V_UNCONNECTED_5201, SV2V_UNCONNECTED_5202, SV2V_UNCONNECTED_5203, SV2V_UNCONNECTED_5204, SV2V_UNCONNECTED_5205, SV2V_UNCONNECTED_5206, SV2V_UNCONNECTED_5207, SV2V_UNCONNECTED_5208, SV2V_UNCONNECTED_5209, SV2V_UNCONNECTED_5210, SV2V_UNCONNECTED_5211, SV2V_UNCONNECTED_5212, SV2V_UNCONNECTED_5213, SV2V_UNCONNECTED_5214, SV2V_UNCONNECTED_5215, SV2V_UNCONNECTED_5216, SV2V_UNCONNECTED_5217, SV2V_UNCONNECTED_5218, SV2V_UNCONNECTED_5219, SV2V_UNCONNECTED_5220, SV2V_UNCONNECTED_5221, SV2V_UNCONNECTED_5222, SV2V_UNCONNECTED_5223, SV2V_UNCONNECTED_5224, SV2V_UNCONNECTED_5225, SV2V_UNCONNECTED_5226, SV2V_UNCONNECTED_5227, SV2V_UNCONNECTED_5228, SV2V_UNCONNECTED_5229, SV2V_UNCONNECTED_5230, SV2V_UNCONNECTED_5231, SV2V_UNCONNECTED_5232, SV2V_UNCONNECTED_5233, SV2V_UNCONNECTED_5234, SV2V_UNCONNECTED_5235, SV2V_UNCONNECTED_5236, SV2V_UNCONNECTED_5237, SV2V_UNCONNECTED_5238, SV2V_UNCONNECTED_5239, SV2V_UNCONNECTED_5240, SV2V_UNCONNECTED_5241, SV2V_UNCONNECTED_5242, SV2V_UNCONNECTED_5243, SV2V_UNCONNECTED_5244, SV2V_UNCONNECTED_5245, SV2V_UNCONNECTED_5246, SV2V_UNCONNECTED_5247, SV2V_UNCONNECTED_5248, SV2V_UNCONNECTED_5249, SV2V_UNCONNECTED_5250, SV2V_UNCONNECTED_5251, SV2V_UNCONNECTED_5252, SV2V_UNCONNECTED_5253, SV2V_UNCONNECTED_5254, SV2V_UNCONNECTED_5255, SV2V_UNCONNECTED_5256, SV2V_UNCONNECTED_5257, SV2V_UNCONNECTED_5258, SV2V_UNCONNECTED_5259, SV2V_UNCONNECTED_5260, SV2V_UNCONNECTED_5261, SV2V_UNCONNECTED_5262, SV2V_UNCONNECTED_5263, SV2V_UNCONNECTED_5264, SV2V_UNCONNECTED_5265, SV2V_UNCONNECTED_5266, SV2V_UNCONNECTED_5267, SV2V_UNCONNECTED_5268, SV2V_UNCONNECTED_5269, SV2V_UNCONNECTED_5270, SV2V_UNCONNECTED_5271, SV2V_UNCONNECTED_5272, SV2V_UNCONNECTED_5273, SV2V_UNCONNECTED_5274, SV2V_UNCONNECTED_5275, SV2V_UNCONNECTED_5276, SV2V_UNCONNECTED_5277, SV2V_UNCONNECTED_5278, SV2V_UNCONNECTED_5279, SV2V_UNCONNECTED_5280, SV2V_UNCONNECTED_5281, SV2V_UNCONNECTED_5282, SV2V_UNCONNECTED_5283, SV2V_UNCONNECTED_5284, SV2V_UNCONNECTED_5285, SV2V_UNCONNECTED_5286, SV2V_UNCONNECTED_5287, SV2V_UNCONNECTED_5288, SV2V_UNCONNECTED_5289, SV2V_UNCONNECTED_5290, SV2V_UNCONNECTED_5291, SV2V_UNCONNECTED_5292, SV2V_UNCONNECTED_5293, SV2V_UNCONNECTED_5294, SV2V_UNCONNECTED_5295, SV2V_UNCONNECTED_5296, SV2V_UNCONNECTED_5297, SV2V_UNCONNECTED_5298, SV2V_UNCONNECTED_5299, SV2V_UNCONNECTED_5300, SV2V_UNCONNECTED_5301, SV2V_UNCONNECTED_5302, SV2V_UNCONNECTED_5303, SV2V_UNCONNECTED_5304, SV2V_UNCONNECTED_5305, SV2V_UNCONNECTED_5306, SV2V_UNCONNECTED_5307, SV2V_UNCONNECTED_5308, SV2V_UNCONNECTED_5309, SV2V_UNCONNECTED_5310, SV2V_UNCONNECTED_5311, SV2V_UNCONNECTED_5312, SV2V_UNCONNECTED_5313, SV2V_UNCONNECTED_5314, SV2V_UNCONNECTED_5315, SV2V_UNCONNECTED_5316, SV2V_UNCONNECTED_5317, SV2V_UNCONNECTED_5318, SV2V_UNCONNECTED_5319, SV2V_UNCONNECTED_5320, SV2V_UNCONNECTED_5321, SV2V_UNCONNECTED_5322, SV2V_UNCONNECTED_5323, SV2V_UNCONNECTED_5324, SV2V_UNCONNECTED_5325, SV2V_UNCONNECTED_5326, SV2V_UNCONNECTED_5327, SV2V_UNCONNECTED_5328, SV2V_UNCONNECTED_5329, SV2V_UNCONNECTED_5330, SV2V_UNCONNECTED_5331, SV2V_UNCONNECTED_5332, SV2V_UNCONNECTED_5333, SV2V_UNCONNECTED_5334, SV2V_UNCONNECTED_5335, SV2V_UNCONNECTED_5336, SV2V_UNCONNECTED_5337, SV2V_UNCONNECTED_5338, SV2V_UNCONNECTED_5339, SV2V_UNCONNECTED_5340, SV2V_UNCONNECTED_5341, SV2V_UNCONNECTED_5342, SV2V_UNCONNECTED_5343, SV2V_UNCONNECTED_5344, SV2V_UNCONNECTED_5345, SV2V_UNCONNECTED_5346, SV2V_UNCONNECTED_5347, SV2V_UNCONNECTED_5348, SV2V_UNCONNECTED_5349, SV2V_UNCONNECTED_5350, SV2V_UNCONNECTED_5351, SV2V_UNCONNECTED_5352, SV2V_UNCONNECTED_5353, SV2V_UNCONNECTED_5354, SV2V_UNCONNECTED_5355, SV2V_UNCONNECTED_5356, SV2V_UNCONNECTED_5357, SV2V_UNCONNECTED_5358, SV2V_UNCONNECTED_5359, SV2V_UNCONNECTED_5360, SV2V_UNCONNECTED_5361, SV2V_UNCONNECTED_5362, SV2V_UNCONNECTED_5363, SV2V_UNCONNECTED_5364, SV2V_UNCONNECTED_5365, SV2V_UNCONNECTED_5366, SV2V_UNCONNECTED_5367, SV2V_UNCONNECTED_5368, SV2V_UNCONNECTED_5369, SV2V_UNCONNECTED_5370, SV2V_UNCONNECTED_5371, SV2V_UNCONNECTED_5372, SV2V_UNCONNECTED_5373, SV2V_UNCONNECTED_5374, SV2V_UNCONNECTED_5375, SV2V_UNCONNECTED_5376, SV2V_UNCONNECTED_5377, SV2V_UNCONNECTED_5378, SV2V_UNCONNECTED_5379, SV2V_UNCONNECTED_5380, SV2V_UNCONNECTED_5381, SV2V_UNCONNECTED_5382, SV2V_UNCONNECTED_5383, SV2V_UNCONNECTED_5384, SV2V_UNCONNECTED_5385, SV2V_UNCONNECTED_5386, SV2V_UNCONNECTED_5387, SV2V_UNCONNECTED_5388, SV2V_UNCONNECTED_5389, SV2V_UNCONNECTED_5390, SV2V_UNCONNECTED_5391, SV2V_UNCONNECTED_5392, SV2V_UNCONNECTED_5393, SV2V_UNCONNECTED_5394, SV2V_UNCONNECTED_5395, SV2V_UNCONNECTED_5396, SV2V_UNCONNECTED_5397, SV2V_UNCONNECTED_5398, SV2V_UNCONNECTED_5399, SV2V_UNCONNECTED_5400, SV2V_UNCONNECTED_5401, SV2V_UNCONNECTED_5402, SV2V_UNCONNECTED_5403, SV2V_UNCONNECTED_5404, SV2V_UNCONNECTED_5405, SV2V_UNCONNECTED_5406, SV2V_UNCONNECTED_5407, SV2V_UNCONNECTED_5408, SV2V_UNCONNECTED_5409, SV2V_UNCONNECTED_5410, SV2V_UNCONNECTED_5411, SV2V_UNCONNECTED_5412, SV2V_UNCONNECTED_5413, SV2V_UNCONNECTED_5414, SV2V_UNCONNECTED_5415, SV2V_UNCONNECTED_5416, SV2V_UNCONNECTED_5417, SV2V_UNCONNECTED_5418, SV2V_UNCONNECTED_5419, SV2V_UNCONNECTED_5420, SV2V_UNCONNECTED_5421, SV2V_UNCONNECTED_5422, SV2V_UNCONNECTED_5423, SV2V_UNCONNECTED_5424, SV2V_UNCONNECTED_5425, SV2V_UNCONNECTED_5426, SV2V_UNCONNECTED_5427, SV2V_UNCONNECTED_5428, SV2V_UNCONNECTED_5429, SV2V_UNCONNECTED_5430, SV2V_UNCONNECTED_5431, SV2V_UNCONNECTED_5432, SV2V_UNCONNECTED_5433, SV2V_UNCONNECTED_5434, SV2V_UNCONNECTED_5435, SV2V_UNCONNECTED_5436, SV2V_UNCONNECTED_5437, SV2V_UNCONNECTED_5438, SV2V_UNCONNECTED_5439, SV2V_UNCONNECTED_5440, SV2V_UNCONNECTED_5441, SV2V_UNCONNECTED_5442, SV2V_UNCONNECTED_5443, SV2V_UNCONNECTED_5444, SV2V_UNCONNECTED_5445, SV2V_UNCONNECTED_5446, SV2V_UNCONNECTED_5447, SV2V_UNCONNECTED_5448, SV2V_UNCONNECTED_5449, SV2V_UNCONNECTED_5450, SV2V_UNCONNECTED_5451, SV2V_UNCONNECTED_5452, SV2V_UNCONNECTED_5453, SV2V_UNCONNECTED_5454, SV2V_UNCONNECTED_5455, SV2V_UNCONNECTED_5456, SV2V_UNCONNECTED_5457, SV2V_UNCONNECTED_5458, SV2V_UNCONNECTED_5459, SV2V_UNCONNECTED_5460, SV2V_UNCONNECTED_5461, SV2V_UNCONNECTED_5462, SV2V_UNCONNECTED_5463, SV2V_UNCONNECTED_5464, SV2V_UNCONNECTED_5465, SV2V_UNCONNECTED_5466, SV2V_UNCONNECTED_5467, SV2V_UNCONNECTED_5468, SV2V_UNCONNECTED_5469, SV2V_UNCONNECTED_5470, SV2V_UNCONNECTED_5471, SV2V_UNCONNECTED_5472, SV2V_UNCONNECTED_5473, SV2V_UNCONNECTED_5474, SV2V_UNCONNECTED_5475, SV2V_UNCONNECTED_5476, SV2V_UNCONNECTED_5477, SV2V_UNCONNECTED_5478, SV2V_UNCONNECTED_5479, SV2V_UNCONNECTED_5480, SV2V_UNCONNECTED_5481, SV2V_UNCONNECTED_5482, SV2V_UNCONNECTED_5483, SV2V_UNCONNECTED_5484, SV2V_UNCONNECTED_5485, SV2V_UNCONNECTED_5486, SV2V_UNCONNECTED_5487, SV2V_UNCONNECTED_5488, SV2V_UNCONNECTED_5489, SV2V_UNCONNECTED_5490, SV2V_UNCONNECTED_5491, SV2V_UNCONNECTED_5492, SV2V_UNCONNECTED_5493, SV2V_UNCONNECTED_5494, SV2V_UNCONNECTED_5495, SV2V_UNCONNECTED_5496, SV2V_UNCONNECTED_5497, SV2V_UNCONNECTED_5498, SV2V_UNCONNECTED_5499, SV2V_UNCONNECTED_5500, SV2V_UNCONNECTED_5501, SV2V_UNCONNECTED_5502, SV2V_UNCONNECTED_5503, SV2V_UNCONNECTED_5504, SV2V_UNCONNECTED_5505, SV2V_UNCONNECTED_5506, SV2V_UNCONNECTED_5507, SV2V_UNCONNECTED_5508, SV2V_UNCONNECTED_5509, SV2V_UNCONNECTED_5510, SV2V_UNCONNECTED_5511, SV2V_UNCONNECTED_5512, SV2V_UNCONNECTED_5513, SV2V_UNCONNECTED_5514, SV2V_UNCONNECTED_5515, SV2V_UNCONNECTED_5516, SV2V_UNCONNECTED_5517, SV2V_UNCONNECTED_5518, SV2V_UNCONNECTED_5519, SV2V_UNCONNECTED_5520, SV2V_UNCONNECTED_5521, SV2V_UNCONNECTED_5522, SV2V_UNCONNECTED_5523, SV2V_UNCONNECTED_5524, SV2V_UNCONNECTED_5525, SV2V_UNCONNECTED_5526, SV2V_UNCONNECTED_5527, SV2V_UNCONNECTED_5528, SV2V_UNCONNECTED_5529, SV2V_UNCONNECTED_5530, SV2V_UNCONNECTED_5531, SV2V_UNCONNECTED_5532, SV2V_UNCONNECTED_5533, SV2V_UNCONNECTED_5534, SV2V_UNCONNECTED_5535, SV2V_UNCONNECTED_5536, SV2V_UNCONNECTED_5537, SV2V_UNCONNECTED_5538, SV2V_UNCONNECTED_5539, SV2V_UNCONNECTED_5540, SV2V_UNCONNECTED_5541, SV2V_UNCONNECTED_5542, SV2V_UNCONNECTED_5543, SV2V_UNCONNECTED_5544, SV2V_UNCONNECTED_5545, SV2V_UNCONNECTED_5546, SV2V_UNCONNECTED_5547, SV2V_UNCONNECTED_5548, SV2V_UNCONNECTED_5549, SV2V_UNCONNECTED_5550, SV2V_UNCONNECTED_5551, SV2V_UNCONNECTED_5552, SV2V_UNCONNECTED_5553, SV2V_UNCONNECTED_5554, SV2V_UNCONNECTED_5555, SV2V_UNCONNECTED_5556, SV2V_UNCONNECTED_5557, SV2V_UNCONNECTED_5558, SV2V_UNCONNECTED_5559, SV2V_UNCONNECTED_5560, SV2V_UNCONNECTED_5561, SV2V_UNCONNECTED_5562, SV2V_UNCONNECTED_5563, SV2V_UNCONNECTED_5564, SV2V_UNCONNECTED_5565, SV2V_UNCONNECTED_5566, SV2V_UNCONNECTED_5567, SV2V_UNCONNECTED_5568, SV2V_UNCONNECTED_5569, SV2V_UNCONNECTED_5570, SV2V_UNCONNECTED_5571, SV2V_UNCONNECTED_5572, SV2V_UNCONNECTED_5573, SV2V_UNCONNECTED_5574, SV2V_UNCONNECTED_5575, SV2V_UNCONNECTED_5576, SV2V_UNCONNECTED_5577, SV2V_UNCONNECTED_5578, SV2V_UNCONNECTED_5579, SV2V_UNCONNECTED_5580, SV2V_UNCONNECTED_5581, SV2V_UNCONNECTED_5582, SV2V_UNCONNECTED_5583, SV2V_UNCONNECTED_5584, SV2V_UNCONNECTED_5585, SV2V_UNCONNECTED_5586, SV2V_UNCONNECTED_5587, SV2V_UNCONNECTED_5588, SV2V_UNCONNECTED_5589, SV2V_UNCONNECTED_5590, SV2V_UNCONNECTED_5591, SV2V_UNCONNECTED_5592, SV2V_UNCONNECTED_5593, SV2V_UNCONNECTED_5594, SV2V_UNCONNECTED_5595, SV2V_UNCONNECTED_5596, SV2V_UNCONNECTED_5597, SV2V_UNCONNECTED_5598, SV2V_UNCONNECTED_5599, SV2V_UNCONNECTED_5600, SV2V_UNCONNECTED_5601, SV2V_UNCONNECTED_5602, SV2V_UNCONNECTED_5603, SV2V_UNCONNECTED_5604, SV2V_UNCONNECTED_5605, SV2V_UNCONNECTED_5606, SV2V_UNCONNECTED_5607, SV2V_UNCONNECTED_5608, SV2V_UNCONNECTED_5609, SV2V_UNCONNECTED_5610, SV2V_UNCONNECTED_5611, SV2V_UNCONNECTED_5612, SV2V_UNCONNECTED_5613, SV2V_UNCONNECTED_5614, SV2V_UNCONNECTED_5615, SV2V_UNCONNECTED_5616, SV2V_UNCONNECTED_5617, SV2V_UNCONNECTED_5618, SV2V_UNCONNECTED_5619, SV2V_UNCONNECTED_5620, SV2V_UNCONNECTED_5621, SV2V_UNCONNECTED_5622, SV2V_UNCONNECTED_5623, SV2V_UNCONNECTED_5624, SV2V_UNCONNECTED_5625, SV2V_UNCONNECTED_5626, SV2V_UNCONNECTED_5627, SV2V_UNCONNECTED_5628, SV2V_UNCONNECTED_5629, SV2V_UNCONNECTED_5630, SV2V_UNCONNECTED_5631, SV2V_UNCONNECTED_5632, SV2V_UNCONNECTED_5633, SV2V_UNCONNECTED_5634, SV2V_UNCONNECTED_5635, SV2V_UNCONNECTED_5636, SV2V_UNCONNECTED_5637, SV2V_UNCONNECTED_5638, SV2V_UNCONNECTED_5639, SV2V_UNCONNECTED_5640, SV2V_UNCONNECTED_5641, SV2V_UNCONNECTED_5642, SV2V_UNCONNECTED_5643, SV2V_UNCONNECTED_5644, SV2V_UNCONNECTED_5645, SV2V_UNCONNECTED_5646, SV2V_UNCONNECTED_5647, SV2V_UNCONNECTED_5648, SV2V_UNCONNECTED_5649, SV2V_UNCONNECTED_5650, SV2V_UNCONNECTED_5651, SV2V_UNCONNECTED_5652, SV2V_UNCONNECTED_5653, SV2V_UNCONNECTED_5654, SV2V_UNCONNECTED_5655, SV2V_UNCONNECTED_5656, SV2V_UNCONNECTED_5657, SV2V_UNCONNECTED_5658, SV2V_UNCONNECTED_5659, SV2V_UNCONNECTED_5660, SV2V_UNCONNECTED_5661, SV2V_UNCONNECTED_5662, SV2V_UNCONNECTED_5663, SV2V_UNCONNECTED_5664, SV2V_UNCONNECTED_5665, SV2V_UNCONNECTED_5666, SV2V_UNCONNECTED_5667, SV2V_UNCONNECTED_5668, SV2V_UNCONNECTED_5669, SV2V_UNCONNECTED_5670, SV2V_UNCONNECTED_5671, SV2V_UNCONNECTED_5672, SV2V_UNCONNECTED_5673, SV2V_UNCONNECTED_5674, SV2V_UNCONNECTED_5675, SV2V_UNCONNECTED_5676, SV2V_UNCONNECTED_5677, SV2V_UNCONNECTED_5678, SV2V_UNCONNECTED_5679, SV2V_UNCONNECTED_5680, SV2V_UNCONNECTED_5681, SV2V_UNCONNECTED_5682, SV2V_UNCONNECTED_5683, SV2V_UNCONNECTED_5684, SV2V_UNCONNECTED_5685, SV2V_UNCONNECTED_5686, SV2V_UNCONNECTED_5687, SV2V_UNCONNECTED_5688, SV2V_UNCONNECTED_5689, SV2V_UNCONNECTED_5690, SV2V_UNCONNECTED_5691, SV2V_UNCONNECTED_5692, SV2V_UNCONNECTED_5693, SV2V_UNCONNECTED_5694, SV2V_UNCONNECTED_5695, SV2V_UNCONNECTED_5696, SV2V_UNCONNECTED_5697, SV2V_UNCONNECTED_5698, SV2V_UNCONNECTED_5699, SV2V_UNCONNECTED_5700, SV2V_UNCONNECTED_5701, SV2V_UNCONNECTED_5702, SV2V_UNCONNECTED_5703, SV2V_UNCONNECTED_5704, SV2V_UNCONNECTED_5705, SV2V_UNCONNECTED_5706, SV2V_UNCONNECTED_5707, SV2V_UNCONNECTED_5708, SV2V_UNCONNECTED_5709, SV2V_UNCONNECTED_5710, SV2V_UNCONNECTED_5711, SV2V_UNCONNECTED_5712, SV2V_UNCONNECTED_5713, SV2V_UNCONNECTED_5714, SV2V_UNCONNECTED_5715, SV2V_UNCONNECTED_5716, SV2V_UNCONNECTED_5717, SV2V_UNCONNECTED_5718, SV2V_UNCONNECTED_5719, SV2V_UNCONNECTED_5720, SV2V_UNCONNECTED_5721, SV2V_UNCONNECTED_5722, SV2V_UNCONNECTED_5723, SV2V_UNCONNECTED_5724, SV2V_UNCONNECTED_5725, SV2V_UNCONNECTED_5726, SV2V_UNCONNECTED_5727, SV2V_UNCONNECTED_5728, SV2V_UNCONNECTED_5729, SV2V_UNCONNECTED_5730, SV2V_UNCONNECTED_5731, SV2V_UNCONNECTED_5732, SV2V_UNCONNECTED_5733, SV2V_UNCONNECTED_5734, SV2V_UNCONNECTED_5735, SV2V_UNCONNECTED_5736, SV2V_UNCONNECTED_5737, SV2V_UNCONNECTED_5738, SV2V_UNCONNECTED_5739, SV2V_UNCONNECTED_5740, SV2V_UNCONNECTED_5741, SV2V_UNCONNECTED_5742, SV2V_UNCONNECTED_5743, SV2V_UNCONNECTED_5744, SV2V_UNCONNECTED_5745, SV2V_UNCONNECTED_5746, SV2V_UNCONNECTED_5747, SV2V_UNCONNECTED_5748, SV2V_UNCONNECTED_5749, SV2V_UNCONNECTED_5750, SV2V_UNCONNECTED_5751, SV2V_UNCONNECTED_5752, SV2V_UNCONNECTED_5753, SV2V_UNCONNECTED_5754, SV2V_UNCONNECTED_5755, SV2V_UNCONNECTED_5756, SV2V_UNCONNECTED_5757, SV2V_UNCONNECTED_5758, SV2V_UNCONNECTED_5759, SV2V_UNCONNECTED_5760, SV2V_UNCONNECTED_5761, SV2V_UNCONNECTED_5762, SV2V_UNCONNECTED_5763, SV2V_UNCONNECTED_5764, SV2V_UNCONNECTED_5765, SV2V_UNCONNECTED_5766, SV2V_UNCONNECTED_5767, SV2V_UNCONNECTED_5768, SV2V_UNCONNECTED_5769, SV2V_UNCONNECTED_5770, SV2V_UNCONNECTED_5771, SV2V_UNCONNECTED_5772, SV2V_UNCONNECTED_5773, SV2V_UNCONNECTED_5774, SV2V_UNCONNECTED_5775, SV2V_UNCONNECTED_5776, SV2V_UNCONNECTED_5777, SV2V_UNCONNECTED_5778, SV2V_UNCONNECTED_5779, SV2V_UNCONNECTED_5780, SV2V_UNCONNECTED_5781, SV2V_UNCONNECTED_5782, SV2V_UNCONNECTED_5783, SV2V_UNCONNECTED_5784, SV2V_UNCONNECTED_5785, SV2V_UNCONNECTED_5786, SV2V_UNCONNECTED_5787, SV2V_UNCONNECTED_5788, SV2V_UNCONNECTED_5789, SV2V_UNCONNECTED_5790, SV2V_UNCONNECTED_5791, SV2V_UNCONNECTED_5792, SV2V_UNCONNECTED_5793, SV2V_UNCONNECTED_5794, SV2V_UNCONNECTED_5795, SV2V_UNCONNECTED_5796, SV2V_UNCONNECTED_5797, SV2V_UNCONNECTED_5798, SV2V_UNCONNECTED_5799, SV2V_UNCONNECTED_5800, SV2V_UNCONNECTED_5801, SV2V_UNCONNECTED_5802, SV2V_UNCONNECTED_5803, SV2V_UNCONNECTED_5804, SV2V_UNCONNECTED_5805, SV2V_UNCONNECTED_5806, SV2V_UNCONNECTED_5807, SV2V_UNCONNECTED_5808, SV2V_UNCONNECTED_5809, SV2V_UNCONNECTED_5810, SV2V_UNCONNECTED_5811, SV2V_UNCONNECTED_5812, SV2V_UNCONNECTED_5813, SV2V_UNCONNECTED_5814, SV2V_UNCONNECTED_5815, SV2V_UNCONNECTED_5816, SV2V_UNCONNECTED_5817, SV2V_UNCONNECTED_5818, SV2V_UNCONNECTED_5819, SV2V_UNCONNECTED_5820, SV2V_UNCONNECTED_5821, SV2V_UNCONNECTED_5822, SV2V_UNCONNECTED_5823, SV2V_UNCONNECTED_5824, SV2V_UNCONNECTED_5825, SV2V_UNCONNECTED_5826, SV2V_UNCONNECTED_5827, SV2V_UNCONNECTED_5828, SV2V_UNCONNECTED_5829, SV2V_UNCONNECTED_5830, SV2V_UNCONNECTED_5831, SV2V_UNCONNECTED_5832, SV2V_UNCONNECTED_5833, SV2V_UNCONNECTED_5834, SV2V_UNCONNECTED_5835, SV2V_UNCONNECTED_5836, SV2V_UNCONNECTED_5837, SV2V_UNCONNECTED_5838, SV2V_UNCONNECTED_5839, SV2V_UNCONNECTED_5840, SV2V_UNCONNECTED_5841, SV2V_UNCONNECTED_5842, SV2V_UNCONNECTED_5843, SV2V_UNCONNECTED_5844, SV2V_UNCONNECTED_5845, SV2V_UNCONNECTED_5846, SV2V_UNCONNECTED_5847, SV2V_UNCONNECTED_5848, SV2V_UNCONNECTED_5849, SV2V_UNCONNECTED_5850, SV2V_UNCONNECTED_5851, SV2V_UNCONNECTED_5852, SV2V_UNCONNECTED_5853, SV2V_UNCONNECTED_5854, SV2V_UNCONNECTED_5855, SV2V_UNCONNECTED_5856, SV2V_UNCONNECTED_5857, SV2V_UNCONNECTED_5858, SV2V_UNCONNECTED_5859, SV2V_UNCONNECTED_5860, SV2V_UNCONNECTED_5861, SV2V_UNCONNECTED_5862, SV2V_UNCONNECTED_5863, SV2V_UNCONNECTED_5864, SV2V_UNCONNECTED_5865, SV2V_UNCONNECTED_5866, SV2V_UNCONNECTED_5867, SV2V_UNCONNECTED_5868, SV2V_UNCONNECTED_5869, SV2V_UNCONNECTED_5870, SV2V_UNCONNECTED_5871, SV2V_UNCONNECTED_5872, SV2V_UNCONNECTED_5873, SV2V_UNCONNECTED_5874, SV2V_UNCONNECTED_5875, SV2V_UNCONNECTED_5876, SV2V_UNCONNECTED_5877, SV2V_UNCONNECTED_5878, SV2V_UNCONNECTED_5879, SV2V_UNCONNECTED_5880, SV2V_UNCONNECTED_5881, SV2V_UNCONNECTED_5882, SV2V_UNCONNECTED_5883, SV2V_UNCONNECTED_5884, SV2V_UNCONNECTED_5885, SV2V_UNCONNECTED_5886, SV2V_UNCONNECTED_5887, SV2V_UNCONNECTED_5888, SV2V_UNCONNECTED_5889, SV2V_UNCONNECTED_5890, SV2V_UNCONNECTED_5891, SV2V_UNCONNECTED_5892, SV2V_UNCONNECTED_5893, SV2V_UNCONNECTED_5894, SV2V_UNCONNECTED_5895, SV2V_UNCONNECTED_5896, SV2V_UNCONNECTED_5897, SV2V_UNCONNECTED_5898, SV2V_UNCONNECTED_5899, SV2V_UNCONNECTED_5900, SV2V_UNCONNECTED_5901, SV2V_UNCONNECTED_5902, SV2V_UNCONNECTED_5903, SV2V_UNCONNECTED_5904, SV2V_UNCONNECTED_5905, SV2V_UNCONNECTED_5906, SV2V_UNCONNECTED_5907, SV2V_UNCONNECTED_5908, SV2V_UNCONNECTED_5909, SV2V_UNCONNECTED_5910, SV2V_UNCONNECTED_5911, SV2V_UNCONNECTED_5912, SV2V_UNCONNECTED_5913, SV2V_UNCONNECTED_5914, SV2V_UNCONNECTED_5915, SV2V_UNCONNECTED_5916, SV2V_UNCONNECTED_5917, SV2V_UNCONNECTED_5918, SV2V_UNCONNECTED_5919, SV2V_UNCONNECTED_5920, SV2V_UNCONNECTED_5921, SV2V_UNCONNECTED_5922, SV2V_UNCONNECTED_5923, SV2V_UNCONNECTED_5924, SV2V_UNCONNECTED_5925, SV2V_UNCONNECTED_5926, SV2V_UNCONNECTED_5927, SV2V_UNCONNECTED_5928, SV2V_UNCONNECTED_5929, SV2V_UNCONNECTED_5930, SV2V_UNCONNECTED_5931, SV2V_UNCONNECTED_5932, SV2V_UNCONNECTED_5933, SV2V_UNCONNECTED_5934, SV2V_UNCONNECTED_5935, SV2V_UNCONNECTED_5936, SV2V_UNCONNECTED_5937, SV2V_UNCONNECTED_5938, SV2V_UNCONNECTED_5939, SV2V_UNCONNECTED_5940, SV2V_UNCONNECTED_5941, SV2V_UNCONNECTED_5942, SV2V_UNCONNECTED_5943, SV2V_UNCONNECTED_5944, SV2V_UNCONNECTED_5945, SV2V_UNCONNECTED_5946, SV2V_UNCONNECTED_5947, SV2V_UNCONNECTED_5948, SV2V_UNCONNECTED_5949, SV2V_UNCONNECTED_5950, SV2V_UNCONNECTED_5951, SV2V_UNCONNECTED_5952, SV2V_UNCONNECTED_5953, SV2V_UNCONNECTED_5954, SV2V_UNCONNECTED_5955, SV2V_UNCONNECTED_5956, SV2V_UNCONNECTED_5957, SV2V_UNCONNECTED_5958, SV2V_UNCONNECTED_5959, SV2V_UNCONNECTED_5960, SV2V_UNCONNECTED_5961, SV2V_UNCONNECTED_5962, SV2V_UNCONNECTED_5963, SV2V_UNCONNECTED_5964, SV2V_UNCONNECTED_5965, SV2V_UNCONNECTED_5966, SV2V_UNCONNECTED_5967, SV2V_UNCONNECTED_5968, SV2V_UNCONNECTED_5969, SV2V_UNCONNECTED_5970, SV2V_UNCONNECTED_5971, SV2V_UNCONNECTED_5972, SV2V_UNCONNECTED_5973, SV2V_UNCONNECTED_5974, SV2V_UNCONNECTED_5975, SV2V_UNCONNECTED_5976, SV2V_UNCONNECTED_5977, SV2V_UNCONNECTED_5978, SV2V_UNCONNECTED_5979, SV2V_UNCONNECTED_5980, SV2V_UNCONNECTED_5981, SV2V_UNCONNECTED_5982, SV2V_UNCONNECTED_5983, SV2V_UNCONNECTED_5984, SV2V_UNCONNECTED_5985, SV2V_UNCONNECTED_5986, SV2V_UNCONNECTED_5987, SV2V_UNCONNECTED_5988, SV2V_UNCONNECTED_5989, SV2V_UNCONNECTED_5990, SV2V_UNCONNECTED_5991, SV2V_UNCONNECTED_5992, SV2V_UNCONNECTED_5993, SV2V_UNCONNECTED_5994, SV2V_UNCONNECTED_5995, SV2V_UNCONNECTED_5996, SV2V_UNCONNECTED_5997, SV2V_UNCONNECTED_5998, SV2V_UNCONNECTED_5999, SV2V_UNCONNECTED_6000, SV2V_UNCONNECTED_6001, SV2V_UNCONNECTED_6002, SV2V_UNCONNECTED_6003, SV2V_UNCONNECTED_6004, SV2V_UNCONNECTED_6005, SV2V_UNCONNECTED_6006, SV2V_UNCONNECTED_6007, SV2V_UNCONNECTED_6008, SV2V_UNCONNECTED_6009, SV2V_UNCONNECTED_6010, SV2V_UNCONNECTED_6011, SV2V_UNCONNECTED_6012, SV2V_UNCONNECTED_6013, SV2V_UNCONNECTED_6014, SV2V_UNCONNECTED_6015, SV2V_UNCONNECTED_6016, SV2V_UNCONNECTED_6017, SV2V_UNCONNECTED_6018, SV2V_UNCONNECTED_6019, SV2V_UNCONNECTED_6020, SV2V_UNCONNECTED_6021, SV2V_UNCONNECTED_6022, SV2V_UNCONNECTED_6023, SV2V_UNCONNECTED_6024, SV2V_UNCONNECTED_6025, SV2V_UNCONNECTED_6026, SV2V_UNCONNECTED_6027, SV2V_UNCONNECTED_6028, SV2V_UNCONNECTED_6029, SV2V_UNCONNECTED_6030, SV2V_UNCONNECTED_6031, SV2V_UNCONNECTED_6032, SV2V_UNCONNECTED_6033, SV2V_UNCONNECTED_6034, SV2V_UNCONNECTED_6035, SV2V_UNCONNECTED_6036, SV2V_UNCONNECTED_6037, SV2V_UNCONNECTED_6038, SV2V_UNCONNECTED_6039, SV2V_UNCONNECTED_6040, SV2V_UNCONNECTED_6041, SV2V_UNCONNECTED_6042, SV2V_UNCONNECTED_6043, SV2V_UNCONNECTED_6044, SV2V_UNCONNECTED_6045, SV2V_UNCONNECTED_6046, SV2V_UNCONNECTED_6047, SV2V_UNCONNECTED_6048, SV2V_UNCONNECTED_6049, SV2V_UNCONNECTED_6050, SV2V_UNCONNECTED_6051, SV2V_UNCONNECTED_6052, SV2V_UNCONNECTED_6053, SV2V_UNCONNECTED_6054, SV2V_UNCONNECTED_6055, SV2V_UNCONNECTED_6056, SV2V_UNCONNECTED_6057, SV2V_UNCONNECTED_6058, SV2V_UNCONNECTED_6059, SV2V_UNCONNECTED_6060, SV2V_UNCONNECTED_6061, SV2V_UNCONNECTED_6062, SV2V_UNCONNECTED_6063, SV2V_UNCONNECTED_6064, SV2V_UNCONNECTED_6065, SV2V_UNCONNECTED_6066, SV2V_UNCONNECTED_6067, SV2V_UNCONNECTED_6068, SV2V_UNCONNECTED_6069, SV2V_UNCONNECTED_6070, SV2V_UNCONNECTED_6071, SV2V_UNCONNECTED_6072, SV2V_UNCONNECTED_6073, SV2V_UNCONNECTED_6074, SV2V_UNCONNECTED_6075, SV2V_UNCONNECTED_6076, SV2V_UNCONNECTED_6077, SV2V_UNCONNECTED_6078, SV2V_UNCONNECTED_6079, SV2V_UNCONNECTED_6080, SV2V_UNCONNECTED_6081, SV2V_UNCONNECTED_6082, SV2V_UNCONNECTED_6083, SV2V_UNCONNECTED_6084, SV2V_UNCONNECTED_6085, SV2V_UNCONNECTED_6086, SV2V_UNCONNECTED_6087, SV2V_UNCONNECTED_6088, SV2V_UNCONNECTED_6089, SV2V_UNCONNECTED_6090, SV2V_UNCONNECTED_6091, SV2V_UNCONNECTED_6092, SV2V_UNCONNECTED_6093, SV2V_UNCONNECTED_6094, SV2V_UNCONNECTED_6095, SV2V_UNCONNECTED_6096, SV2V_UNCONNECTED_6097, SV2V_UNCONNECTED_6098, SV2V_UNCONNECTED_6099, SV2V_UNCONNECTED_6100, SV2V_UNCONNECTED_6101, SV2V_UNCONNECTED_6102, SV2V_UNCONNECTED_6103, SV2V_UNCONNECTED_6104, SV2V_UNCONNECTED_6105, SV2V_UNCONNECTED_6106, SV2V_UNCONNECTED_6107, SV2V_UNCONNECTED_6108, SV2V_UNCONNECTED_6109, SV2V_UNCONNECTED_6110, SV2V_UNCONNECTED_6111, SV2V_UNCONNECTED_6112, SV2V_UNCONNECTED_6113, SV2V_UNCONNECTED_6114, SV2V_UNCONNECTED_6115, SV2V_UNCONNECTED_6116, SV2V_UNCONNECTED_6117, SV2V_UNCONNECTED_6118, SV2V_UNCONNECTED_6119, SV2V_UNCONNECTED_6120, SV2V_UNCONNECTED_6121, SV2V_UNCONNECTED_6122, SV2V_UNCONNECTED_6123, SV2V_UNCONNECTED_6124, SV2V_UNCONNECTED_6125, SV2V_UNCONNECTED_6126, SV2V_UNCONNECTED_6127, SV2V_UNCONNECTED_6128, SV2V_UNCONNECTED_6129, SV2V_UNCONNECTED_6130, SV2V_UNCONNECTED_6131, SV2V_UNCONNECTED_6132, SV2V_UNCONNECTED_6133, SV2V_UNCONNECTED_6134, SV2V_UNCONNECTED_6135, SV2V_UNCONNECTED_6136, SV2V_UNCONNECTED_6137, SV2V_UNCONNECTED_6138, SV2V_UNCONNECTED_6139, SV2V_UNCONNECTED_6140, SV2V_UNCONNECTED_6141, SV2V_UNCONNECTED_6142, SV2V_UNCONNECTED_6143, SV2V_UNCONNECTED_6144, SV2V_UNCONNECTED_6145, SV2V_UNCONNECTED_6146, SV2V_UNCONNECTED_6147, SV2V_UNCONNECTED_6148, SV2V_UNCONNECTED_6149, SV2V_UNCONNECTED_6150, SV2V_UNCONNECTED_6151, SV2V_UNCONNECTED_6152, SV2V_UNCONNECTED_6153, SV2V_UNCONNECTED_6154, SV2V_UNCONNECTED_6155, SV2V_UNCONNECTED_6156, SV2V_UNCONNECTED_6157, SV2V_UNCONNECTED_6158, SV2V_UNCONNECTED_6159, SV2V_UNCONNECTED_6160, SV2V_UNCONNECTED_6161, SV2V_UNCONNECTED_6162, SV2V_UNCONNECTED_6163, SV2V_UNCONNECTED_6164, SV2V_UNCONNECTED_6165, SV2V_UNCONNECTED_6166, SV2V_UNCONNECTED_6167, SV2V_UNCONNECTED_6168, SV2V_UNCONNECTED_6169, SV2V_UNCONNECTED_6170, SV2V_UNCONNECTED_6171, SV2V_UNCONNECTED_6172, SV2V_UNCONNECTED_6173, SV2V_UNCONNECTED_6174, SV2V_UNCONNECTED_6175, SV2V_UNCONNECTED_6176, SV2V_UNCONNECTED_6177, SV2V_UNCONNECTED_6178, SV2V_UNCONNECTED_6179, SV2V_UNCONNECTED_6180, SV2V_UNCONNECTED_6181, SV2V_UNCONNECTED_6182, SV2V_UNCONNECTED_6183, SV2V_UNCONNECTED_6184, SV2V_UNCONNECTED_6185, SV2V_UNCONNECTED_6186, SV2V_UNCONNECTED_6187, SV2V_UNCONNECTED_6188, SV2V_UNCONNECTED_6189, SV2V_UNCONNECTED_6190, SV2V_UNCONNECTED_6191, SV2V_UNCONNECTED_6192, SV2V_UNCONNECTED_6193, SV2V_UNCONNECTED_6194, SV2V_UNCONNECTED_6195, SV2V_UNCONNECTED_6196, SV2V_UNCONNECTED_6197, SV2V_UNCONNECTED_6198, SV2V_UNCONNECTED_6199, SV2V_UNCONNECTED_6200, SV2V_UNCONNECTED_6201, SV2V_UNCONNECTED_6202, SV2V_UNCONNECTED_6203, SV2V_UNCONNECTED_6204, SV2V_UNCONNECTED_6205, SV2V_UNCONNECTED_6206, SV2V_UNCONNECTED_6207, SV2V_UNCONNECTED_6208, SV2V_UNCONNECTED_6209, SV2V_UNCONNECTED_6210, SV2V_UNCONNECTED_6211, SV2V_UNCONNECTED_6212, SV2V_UNCONNECTED_6213, SV2V_UNCONNECTED_6214, SV2V_UNCONNECTED_6215, SV2V_UNCONNECTED_6216, SV2V_UNCONNECTED_6217, SV2V_UNCONNECTED_6218, SV2V_UNCONNECTED_6219, SV2V_UNCONNECTED_6220, SV2V_UNCONNECTED_6221, SV2V_UNCONNECTED_6222, SV2V_UNCONNECTED_6223, SV2V_UNCONNECTED_6224, SV2V_UNCONNECTED_6225, SV2V_UNCONNECTED_6226, SV2V_UNCONNECTED_6227, SV2V_UNCONNECTED_6228, SV2V_UNCONNECTED_6229, SV2V_UNCONNECTED_6230, SV2V_UNCONNECTED_6231, SV2V_UNCONNECTED_6232, SV2V_UNCONNECTED_6233, SV2V_UNCONNECTED_6234, SV2V_UNCONNECTED_6235, SV2V_UNCONNECTED_6236, SV2V_UNCONNECTED_6237, SV2V_UNCONNECTED_6238, SV2V_UNCONNECTED_6239, SV2V_UNCONNECTED_6240, SV2V_UNCONNECTED_6241, SV2V_UNCONNECTED_6242, SV2V_UNCONNECTED_6243, SV2V_UNCONNECTED_6244, SV2V_UNCONNECTED_6245, SV2V_UNCONNECTED_6246, SV2V_UNCONNECTED_6247, SV2V_UNCONNECTED_6248, SV2V_UNCONNECTED_6249, SV2V_UNCONNECTED_6250, SV2V_UNCONNECTED_6251, SV2V_UNCONNECTED_6252, SV2V_UNCONNECTED_6253, SV2V_UNCONNECTED_6254, SV2V_UNCONNECTED_6255, SV2V_UNCONNECTED_6256, SV2V_UNCONNECTED_6257, SV2V_UNCONNECTED_6258, SV2V_UNCONNECTED_6259, SV2V_UNCONNECTED_6260, SV2V_UNCONNECTED_6261, SV2V_UNCONNECTED_6262, SV2V_UNCONNECTED_6263, SV2V_UNCONNECTED_6264, SV2V_UNCONNECTED_6265, SV2V_UNCONNECTED_6266, SV2V_UNCONNECTED_6267, SV2V_UNCONNECTED_6268, SV2V_UNCONNECTED_6269, SV2V_UNCONNECTED_6270, SV2V_UNCONNECTED_6271, SV2V_UNCONNECTED_6272, SV2V_UNCONNECTED_6273, SV2V_UNCONNECTED_6274, SV2V_UNCONNECTED_6275, SV2V_UNCONNECTED_6276, SV2V_UNCONNECTED_6277, SV2V_UNCONNECTED_6278, SV2V_UNCONNECTED_6279, SV2V_UNCONNECTED_6280, SV2V_UNCONNECTED_6281, SV2V_UNCONNECTED_6282, SV2V_UNCONNECTED_6283, SV2V_UNCONNECTED_6284, SV2V_UNCONNECTED_6285, SV2V_UNCONNECTED_6286, SV2V_UNCONNECTED_6287, SV2V_UNCONNECTED_6288, SV2V_UNCONNECTED_6289, SV2V_UNCONNECTED_6290, SV2V_UNCONNECTED_6291, SV2V_UNCONNECTED_6292, SV2V_UNCONNECTED_6293, SV2V_UNCONNECTED_6294, SV2V_UNCONNECTED_6295, SV2V_UNCONNECTED_6296, SV2V_UNCONNECTED_6297, SV2V_UNCONNECTED_6298, SV2V_UNCONNECTED_6299, SV2V_UNCONNECTED_6300, SV2V_UNCONNECTED_6301, SV2V_UNCONNECTED_6302, SV2V_UNCONNECTED_6303, SV2V_UNCONNECTED_6304, SV2V_UNCONNECTED_6305, SV2V_UNCONNECTED_6306, SV2V_UNCONNECTED_6307, SV2V_UNCONNECTED_6308, SV2V_UNCONNECTED_6309, SV2V_UNCONNECTED_6310, SV2V_UNCONNECTED_6311, SV2V_UNCONNECTED_6312, SV2V_UNCONNECTED_6313, SV2V_UNCONNECTED_6314, SV2V_UNCONNECTED_6315, SV2V_UNCONNECTED_6316, SV2V_UNCONNECTED_6317, SV2V_UNCONNECTED_6318, SV2V_UNCONNECTED_6319, SV2V_UNCONNECTED_6320, SV2V_UNCONNECTED_6321, SV2V_UNCONNECTED_6322, SV2V_UNCONNECTED_6323, SV2V_UNCONNECTED_6324, SV2V_UNCONNECTED_6325, SV2V_UNCONNECTED_6326, SV2V_UNCONNECTED_6327, SV2V_UNCONNECTED_6328, SV2V_UNCONNECTED_6329, SV2V_UNCONNECTED_6330, SV2V_UNCONNECTED_6331, SV2V_UNCONNECTED_6332, SV2V_UNCONNECTED_6333, SV2V_UNCONNECTED_6334, SV2V_UNCONNECTED_6335, SV2V_UNCONNECTED_6336, SV2V_UNCONNECTED_6337, SV2V_UNCONNECTED_6338, SV2V_UNCONNECTED_6339, SV2V_UNCONNECTED_6340, SV2V_UNCONNECTED_6341, SV2V_UNCONNECTED_6342, SV2V_UNCONNECTED_6343, SV2V_UNCONNECTED_6344, SV2V_UNCONNECTED_6345, SV2V_UNCONNECTED_6346, SV2V_UNCONNECTED_6347, SV2V_UNCONNECTED_6348, SV2V_UNCONNECTED_6349, SV2V_UNCONNECTED_6350, SV2V_UNCONNECTED_6351, SV2V_UNCONNECTED_6352, SV2V_UNCONNECTED_6353, SV2V_UNCONNECTED_6354, SV2V_UNCONNECTED_6355, SV2V_UNCONNECTED_6356, SV2V_UNCONNECTED_6357, SV2V_UNCONNECTED_6358, SV2V_UNCONNECTED_6359, SV2V_UNCONNECTED_6360, SV2V_UNCONNECTED_6361, SV2V_UNCONNECTED_6362, SV2V_UNCONNECTED_6363, SV2V_UNCONNECTED_6364, SV2V_UNCONNECTED_6365, SV2V_UNCONNECTED_6366, SV2V_UNCONNECTED_6367, SV2V_UNCONNECTED_6368, SV2V_UNCONNECTED_6369, SV2V_UNCONNECTED_6370, SV2V_UNCONNECTED_6371, SV2V_UNCONNECTED_6372, SV2V_UNCONNECTED_6373, SV2V_UNCONNECTED_6374, SV2V_UNCONNECTED_6375, SV2V_UNCONNECTED_6376, SV2V_UNCONNECTED_6377, SV2V_UNCONNECTED_6378, SV2V_UNCONNECTED_6379, SV2V_UNCONNECTED_6380, SV2V_UNCONNECTED_6381, SV2V_UNCONNECTED_6382, SV2V_UNCONNECTED_6383, SV2V_UNCONNECTED_6384, SV2V_UNCONNECTED_6385, SV2V_UNCONNECTED_6386, SV2V_UNCONNECTED_6387, SV2V_UNCONNECTED_6388, SV2V_UNCONNECTED_6389, SV2V_UNCONNECTED_6390, SV2V_UNCONNECTED_6391, SV2V_UNCONNECTED_6392, SV2V_UNCONNECTED_6393, SV2V_UNCONNECTED_6394, SV2V_UNCONNECTED_6395, SV2V_UNCONNECTED_6396, SV2V_UNCONNECTED_6397, SV2V_UNCONNECTED_6398, SV2V_UNCONNECTED_6399, SV2V_UNCONNECTED_6400, SV2V_UNCONNECTED_6401, SV2V_UNCONNECTED_6402, SV2V_UNCONNECTED_6403, SV2V_UNCONNECTED_6404, SV2V_UNCONNECTED_6405, SV2V_UNCONNECTED_6406, SV2V_UNCONNECTED_6407, SV2V_UNCONNECTED_6408, SV2V_UNCONNECTED_6409, SV2V_UNCONNECTED_6410, SV2V_UNCONNECTED_6411, SV2V_UNCONNECTED_6412, SV2V_UNCONNECTED_6413, SV2V_UNCONNECTED_6414, SV2V_UNCONNECTED_6415, SV2V_UNCONNECTED_6416, SV2V_UNCONNECTED_6417, SV2V_UNCONNECTED_6418, SV2V_UNCONNECTED_6419, SV2V_UNCONNECTED_6420, SV2V_UNCONNECTED_6421, SV2V_UNCONNECTED_6422, SV2V_UNCONNECTED_6423, SV2V_UNCONNECTED_6424, SV2V_UNCONNECTED_6425, SV2V_UNCONNECTED_6426, SV2V_UNCONNECTED_6427, SV2V_UNCONNECTED_6428, SV2V_UNCONNECTED_6429, SV2V_UNCONNECTED_6430, SV2V_UNCONNECTED_6431, SV2V_UNCONNECTED_6432, SV2V_UNCONNECTED_6433, SV2V_UNCONNECTED_6434, SV2V_UNCONNECTED_6435, SV2V_UNCONNECTED_6436, SV2V_UNCONNECTED_6437, SV2V_UNCONNECTED_6438, SV2V_UNCONNECTED_6439, SV2V_UNCONNECTED_6440, SV2V_UNCONNECTED_6441, SV2V_UNCONNECTED_6442, SV2V_UNCONNECTED_6443, SV2V_UNCONNECTED_6444, SV2V_UNCONNECTED_6445, SV2V_UNCONNECTED_6446, SV2V_UNCONNECTED_6447, SV2V_UNCONNECTED_6448, SV2V_UNCONNECTED_6449, SV2V_UNCONNECTED_6450, SV2V_UNCONNECTED_6451, SV2V_UNCONNECTED_6452, SV2V_UNCONNECTED_6453, SV2V_UNCONNECTED_6454, SV2V_UNCONNECTED_6455, SV2V_UNCONNECTED_6456, SV2V_UNCONNECTED_6457, SV2V_UNCONNECTED_6458, SV2V_UNCONNECTED_6459, SV2V_UNCONNECTED_6460, SV2V_UNCONNECTED_6461, SV2V_UNCONNECTED_6462, SV2V_UNCONNECTED_6463, SV2V_UNCONNECTED_6464, SV2V_UNCONNECTED_6465, SV2V_UNCONNECTED_6466, SV2V_UNCONNECTED_6467, SV2V_UNCONNECTED_6468, SV2V_UNCONNECTED_6469, SV2V_UNCONNECTED_6470, SV2V_UNCONNECTED_6471, SV2V_UNCONNECTED_6472, SV2V_UNCONNECTED_6473, SV2V_UNCONNECTED_6474, SV2V_UNCONNECTED_6475, SV2V_UNCONNECTED_6476, SV2V_UNCONNECTED_6477, SV2V_UNCONNECTED_6478, SV2V_UNCONNECTED_6479, SV2V_UNCONNECTED_6480, SV2V_UNCONNECTED_6481, SV2V_UNCONNECTED_6482, SV2V_UNCONNECTED_6483, SV2V_UNCONNECTED_6484, SV2V_UNCONNECTED_6485, SV2V_UNCONNECTED_6486, SV2V_UNCONNECTED_6487, SV2V_UNCONNECTED_6488, SV2V_UNCONNECTED_6489, SV2V_UNCONNECTED_6490, SV2V_UNCONNECTED_6491, SV2V_UNCONNECTED_6492, SV2V_UNCONNECTED_6493, SV2V_UNCONNECTED_6494, SV2V_UNCONNECTED_6495, SV2V_UNCONNECTED_6496, SV2V_UNCONNECTED_6497, SV2V_UNCONNECTED_6498, SV2V_UNCONNECTED_6499, SV2V_UNCONNECTED_6500, SV2V_UNCONNECTED_6501, SV2V_UNCONNECTED_6502, SV2V_UNCONNECTED_6503, SV2V_UNCONNECTED_6504, SV2V_UNCONNECTED_6505, SV2V_UNCONNECTED_6506, SV2V_UNCONNECTED_6507, SV2V_UNCONNECTED_6508, SV2V_UNCONNECTED_6509, SV2V_UNCONNECTED_6510, SV2V_UNCONNECTED_6511, SV2V_UNCONNECTED_6512, SV2V_UNCONNECTED_6513, SV2V_UNCONNECTED_6514, SV2V_UNCONNECTED_6515, SV2V_UNCONNECTED_6516, SV2V_UNCONNECTED_6517, SV2V_UNCONNECTED_6518, SV2V_UNCONNECTED_6519, SV2V_UNCONNECTED_6520, SV2V_UNCONNECTED_6521, SV2V_UNCONNECTED_6522, SV2V_UNCONNECTED_6523, SV2V_UNCONNECTED_6524, SV2V_UNCONNECTED_6525, SV2V_UNCONNECTED_6526, SV2V_UNCONNECTED_6527, SV2V_UNCONNECTED_6528, SV2V_UNCONNECTED_6529, SV2V_UNCONNECTED_6530, SV2V_UNCONNECTED_6531, SV2V_UNCONNECTED_6532, SV2V_UNCONNECTED_6533, SV2V_UNCONNECTED_6534, SV2V_UNCONNECTED_6535, SV2V_UNCONNECTED_6536, SV2V_UNCONNECTED_6537, SV2V_UNCONNECTED_6538, SV2V_UNCONNECTED_6539, SV2V_UNCONNECTED_6540, SV2V_UNCONNECTED_6541, SV2V_UNCONNECTED_6542, SV2V_UNCONNECTED_6543, SV2V_UNCONNECTED_6544, SV2V_UNCONNECTED_6545, SV2V_UNCONNECTED_6546, SV2V_UNCONNECTED_6547, SV2V_UNCONNECTED_6548, SV2V_UNCONNECTED_6549, SV2V_UNCONNECTED_6550, SV2V_UNCONNECTED_6551, SV2V_UNCONNECTED_6552, SV2V_UNCONNECTED_6553, SV2V_UNCONNECTED_6554, SV2V_UNCONNECTED_6555, SV2V_UNCONNECTED_6556, SV2V_UNCONNECTED_6557, SV2V_UNCONNECTED_6558, SV2V_UNCONNECTED_6559, SV2V_UNCONNECTED_6560, SV2V_UNCONNECTED_6561, SV2V_UNCONNECTED_6562, SV2V_UNCONNECTED_6563, SV2V_UNCONNECTED_6564, SV2V_UNCONNECTED_6565, SV2V_UNCONNECTED_6566, SV2V_UNCONNECTED_6567, SV2V_UNCONNECTED_6568, SV2V_UNCONNECTED_6569, SV2V_UNCONNECTED_6570, SV2V_UNCONNECTED_6571, SV2V_UNCONNECTED_6572, SV2V_UNCONNECTED_6573, SV2V_UNCONNECTED_6574, SV2V_UNCONNECTED_6575, SV2V_UNCONNECTED_6576, SV2V_UNCONNECTED_6577, SV2V_UNCONNECTED_6578, SV2V_UNCONNECTED_6579, SV2V_UNCONNECTED_6580, SV2V_UNCONNECTED_6581, SV2V_UNCONNECTED_6582, SV2V_UNCONNECTED_6583, SV2V_UNCONNECTED_6584, SV2V_UNCONNECTED_6585, SV2V_UNCONNECTED_6586, SV2V_UNCONNECTED_6587, SV2V_UNCONNECTED_6588, SV2V_UNCONNECTED_6589, SV2V_UNCONNECTED_6590, SV2V_UNCONNECTED_6591, SV2V_UNCONNECTED_6592, SV2V_UNCONNECTED_6593, SV2V_UNCONNECTED_6594, SV2V_UNCONNECTED_6595, SV2V_UNCONNECTED_6596, SV2V_UNCONNECTED_6597, SV2V_UNCONNECTED_6598, SV2V_UNCONNECTED_6599, SV2V_UNCONNECTED_6600, SV2V_UNCONNECTED_6601, SV2V_UNCONNECTED_6602, SV2V_UNCONNECTED_6603, SV2V_UNCONNECTED_6604, SV2V_UNCONNECTED_6605, SV2V_UNCONNECTED_6606, SV2V_UNCONNECTED_6607, SV2V_UNCONNECTED_6608, SV2V_UNCONNECTED_6609, SV2V_UNCONNECTED_6610, SV2V_UNCONNECTED_6611, SV2V_UNCONNECTED_6612, SV2V_UNCONNECTED_6613, SV2V_UNCONNECTED_6614, SV2V_UNCONNECTED_6615, SV2V_UNCONNECTED_6616, SV2V_UNCONNECTED_6617, SV2V_UNCONNECTED_6618, SV2V_UNCONNECTED_6619, SV2V_UNCONNECTED_6620, SV2V_UNCONNECTED_6621, SV2V_UNCONNECTED_6622, SV2V_UNCONNECTED_6623, SV2V_UNCONNECTED_6624, SV2V_UNCONNECTED_6625, SV2V_UNCONNECTED_6626, SV2V_UNCONNECTED_6627, SV2V_UNCONNECTED_6628, SV2V_UNCONNECTED_6629, SV2V_UNCONNECTED_6630, SV2V_UNCONNECTED_6631, SV2V_UNCONNECTED_6632, SV2V_UNCONNECTED_6633, SV2V_UNCONNECTED_6634, SV2V_UNCONNECTED_6635, SV2V_UNCONNECTED_6636, SV2V_UNCONNECTED_6637, SV2V_UNCONNECTED_6638, SV2V_UNCONNECTED_6639, SV2V_UNCONNECTED_6640, SV2V_UNCONNECTED_6641, SV2V_UNCONNECTED_6642, SV2V_UNCONNECTED_6643, SV2V_UNCONNECTED_6644, SV2V_UNCONNECTED_6645, SV2V_UNCONNECTED_6646, SV2V_UNCONNECTED_6647, SV2V_UNCONNECTED_6648, SV2V_UNCONNECTED_6649, SV2V_UNCONNECTED_6650, SV2V_UNCONNECTED_6651, SV2V_UNCONNECTED_6652, SV2V_UNCONNECTED_6653, SV2V_UNCONNECTED_6654, SV2V_UNCONNECTED_6655, SV2V_UNCONNECTED_6656, SV2V_UNCONNECTED_6657, SV2V_UNCONNECTED_6658, SV2V_UNCONNECTED_6659, SV2V_UNCONNECTED_6660, SV2V_UNCONNECTED_6661, SV2V_UNCONNECTED_6662, SV2V_UNCONNECTED_6663, SV2V_UNCONNECTED_6664, SV2V_UNCONNECTED_6665, SV2V_UNCONNECTED_6666, SV2V_UNCONNECTED_6667, SV2V_UNCONNECTED_6668, SV2V_UNCONNECTED_6669, SV2V_UNCONNECTED_6670, SV2V_UNCONNECTED_6671, SV2V_UNCONNECTED_6672, SV2V_UNCONNECTED_6673, SV2V_UNCONNECTED_6674, SV2V_UNCONNECTED_6675, SV2V_UNCONNECTED_6676, SV2V_UNCONNECTED_6677, SV2V_UNCONNECTED_6678, SV2V_UNCONNECTED_6679, SV2V_UNCONNECTED_6680, SV2V_UNCONNECTED_6681, SV2V_UNCONNECTED_6682, SV2V_UNCONNECTED_6683, SV2V_UNCONNECTED_6684, SV2V_UNCONNECTED_6685, SV2V_UNCONNECTED_6686, SV2V_UNCONNECTED_6687, SV2V_UNCONNECTED_6688, SV2V_UNCONNECTED_6689, SV2V_UNCONNECTED_6690, SV2V_UNCONNECTED_6691, SV2V_UNCONNECTED_6692, SV2V_UNCONNECTED_6693, SV2V_UNCONNECTED_6694, SV2V_UNCONNECTED_6695, SV2V_UNCONNECTED_6696, SV2V_UNCONNECTED_6697, SV2V_UNCONNECTED_6698, SV2V_UNCONNECTED_6699, SV2V_UNCONNECTED_6700, SV2V_UNCONNECTED_6701, SV2V_UNCONNECTED_6702, SV2V_UNCONNECTED_6703, SV2V_UNCONNECTED_6704, SV2V_UNCONNECTED_6705, SV2V_UNCONNECTED_6706, SV2V_UNCONNECTED_6707, SV2V_UNCONNECTED_6708, SV2V_UNCONNECTED_6709, SV2V_UNCONNECTED_6710, SV2V_UNCONNECTED_6711, SV2V_UNCONNECTED_6712, SV2V_UNCONNECTED_6713, SV2V_UNCONNECTED_6714, SV2V_UNCONNECTED_6715, SV2V_UNCONNECTED_6716, SV2V_UNCONNECTED_6717, SV2V_UNCONNECTED_6718, SV2V_UNCONNECTED_6719, SV2V_UNCONNECTED_6720, SV2V_UNCONNECTED_6721, SV2V_UNCONNECTED_6722, SV2V_UNCONNECTED_6723, SV2V_UNCONNECTED_6724, SV2V_UNCONNECTED_6725, SV2V_UNCONNECTED_6726, SV2V_UNCONNECTED_6727, SV2V_UNCONNECTED_6728, SV2V_UNCONNECTED_6729, SV2V_UNCONNECTED_6730, SV2V_UNCONNECTED_6731, SV2V_UNCONNECTED_6732, SV2V_UNCONNECTED_6733, SV2V_UNCONNECTED_6734, SV2V_UNCONNECTED_6735, SV2V_UNCONNECTED_6736, SV2V_UNCONNECTED_6737, SV2V_UNCONNECTED_6738, SV2V_UNCONNECTED_6739, SV2V_UNCONNECTED_6740, SV2V_UNCONNECTED_6741, SV2V_UNCONNECTED_6742, SV2V_UNCONNECTED_6743, SV2V_UNCONNECTED_6744, SV2V_UNCONNECTED_6745, SV2V_UNCONNECTED_6746, SV2V_UNCONNECTED_6747, SV2V_UNCONNECTED_6748, SV2V_UNCONNECTED_6749, SV2V_UNCONNECTED_6750, SV2V_UNCONNECTED_6751, SV2V_UNCONNECTED_6752, SV2V_UNCONNECTED_6753, SV2V_UNCONNECTED_6754, SV2V_UNCONNECTED_6755, SV2V_UNCONNECTED_6756, SV2V_UNCONNECTED_6757, SV2V_UNCONNECTED_6758, SV2V_UNCONNECTED_6759, SV2V_UNCONNECTED_6760, SV2V_UNCONNECTED_6761, SV2V_UNCONNECTED_6762, SV2V_UNCONNECTED_6763, SV2V_UNCONNECTED_6764, SV2V_UNCONNECTED_6765, SV2V_UNCONNECTED_6766, SV2V_UNCONNECTED_6767, SV2V_UNCONNECTED_6768, SV2V_UNCONNECTED_6769, SV2V_UNCONNECTED_6770, SV2V_UNCONNECTED_6771, SV2V_UNCONNECTED_6772, SV2V_UNCONNECTED_6773, SV2V_UNCONNECTED_6774, SV2V_UNCONNECTED_6775, SV2V_UNCONNECTED_6776, SV2V_UNCONNECTED_6777, SV2V_UNCONNECTED_6778, SV2V_UNCONNECTED_6779, SV2V_UNCONNECTED_6780, SV2V_UNCONNECTED_6781, SV2V_UNCONNECTED_6782, SV2V_UNCONNECTED_6783, SV2V_UNCONNECTED_6784, SV2V_UNCONNECTED_6785, SV2V_UNCONNECTED_6786, SV2V_UNCONNECTED_6787, SV2V_UNCONNECTED_6788, SV2V_UNCONNECTED_6789, SV2V_UNCONNECTED_6790, SV2V_UNCONNECTED_6791, SV2V_UNCONNECTED_6792, SV2V_UNCONNECTED_6793, SV2V_UNCONNECTED_6794, SV2V_UNCONNECTED_6795, SV2V_UNCONNECTED_6796, SV2V_UNCONNECTED_6797, SV2V_UNCONNECTED_6798, SV2V_UNCONNECTED_6799, SV2V_UNCONNECTED_6800, SV2V_UNCONNECTED_6801, SV2V_UNCONNECTED_6802, SV2V_UNCONNECTED_6803, SV2V_UNCONNECTED_6804, SV2V_UNCONNECTED_6805, SV2V_UNCONNECTED_6806, SV2V_UNCONNECTED_6807, SV2V_UNCONNECTED_6808, SV2V_UNCONNECTED_6809, SV2V_UNCONNECTED_6810, SV2V_UNCONNECTED_6811, SV2V_UNCONNECTED_6812, SV2V_UNCONNECTED_6813, SV2V_UNCONNECTED_6814, SV2V_UNCONNECTED_6815, SV2V_UNCONNECTED_6816, SV2V_UNCONNECTED_6817, SV2V_UNCONNECTED_6818, SV2V_UNCONNECTED_6819, SV2V_UNCONNECTED_6820, SV2V_UNCONNECTED_6821, SV2V_UNCONNECTED_6822, SV2V_UNCONNECTED_6823, SV2V_UNCONNECTED_6824, SV2V_UNCONNECTED_6825, SV2V_UNCONNECTED_6826, SV2V_UNCONNECTED_6827, SV2V_UNCONNECTED_6828, SV2V_UNCONNECTED_6829, SV2V_UNCONNECTED_6830, SV2V_UNCONNECTED_6831, SV2V_UNCONNECTED_6832, SV2V_UNCONNECTED_6833, SV2V_UNCONNECTED_6834, SV2V_UNCONNECTED_6835, SV2V_UNCONNECTED_6836, SV2V_UNCONNECTED_6837, SV2V_UNCONNECTED_6838, SV2V_UNCONNECTED_6839, SV2V_UNCONNECTED_6840, SV2V_UNCONNECTED_6841, SV2V_UNCONNECTED_6842, SV2V_UNCONNECTED_6843, SV2V_UNCONNECTED_6844, SV2V_UNCONNECTED_6845, SV2V_UNCONNECTED_6846, SV2V_UNCONNECTED_6847, SV2V_UNCONNECTED_6848, SV2V_UNCONNECTED_6849, SV2V_UNCONNECTED_6850, SV2V_UNCONNECTED_6851, SV2V_UNCONNECTED_6852, SV2V_UNCONNECTED_6853, SV2V_UNCONNECTED_6854, SV2V_UNCONNECTED_6855, SV2V_UNCONNECTED_6856, SV2V_UNCONNECTED_6857, SV2V_UNCONNECTED_6858, SV2V_UNCONNECTED_6859, SV2V_UNCONNECTED_6860, SV2V_UNCONNECTED_6861, SV2V_UNCONNECTED_6862, SV2V_UNCONNECTED_6863, SV2V_UNCONNECTED_6864, SV2V_UNCONNECTED_6865, SV2V_UNCONNECTED_6866, SV2V_UNCONNECTED_6867, SV2V_UNCONNECTED_6868, SV2V_UNCONNECTED_6869, SV2V_UNCONNECTED_6870, SV2V_UNCONNECTED_6871, SV2V_UNCONNECTED_6872, SV2V_UNCONNECTED_6873, SV2V_UNCONNECTED_6874, SV2V_UNCONNECTED_6875, SV2V_UNCONNECTED_6876, SV2V_UNCONNECTED_6877, SV2V_UNCONNECTED_6878, SV2V_UNCONNECTED_6879, SV2V_UNCONNECTED_6880, SV2V_UNCONNECTED_6881, SV2V_UNCONNECTED_6882, SV2V_UNCONNECTED_6883, SV2V_UNCONNECTED_6884, SV2V_UNCONNECTED_6885, SV2V_UNCONNECTED_6886, SV2V_UNCONNECTED_6887, SV2V_UNCONNECTED_6888, SV2V_UNCONNECTED_6889, SV2V_UNCONNECTED_6890, SV2V_UNCONNECTED_6891, SV2V_UNCONNECTED_6892, SV2V_UNCONNECTED_6893, SV2V_UNCONNECTED_6894, SV2V_UNCONNECTED_6895, SV2V_UNCONNECTED_6896, SV2V_UNCONNECTED_6897, SV2V_UNCONNECTED_6898, SV2V_UNCONNECTED_6899, SV2V_UNCONNECTED_6900, SV2V_UNCONNECTED_6901, SV2V_UNCONNECTED_6902, SV2V_UNCONNECTED_6903, SV2V_UNCONNECTED_6904, SV2V_UNCONNECTED_6905, SV2V_UNCONNECTED_6906, SV2V_UNCONNECTED_6907, SV2V_UNCONNECTED_6908, SV2V_UNCONNECTED_6909, SV2V_UNCONNECTED_6910, SV2V_UNCONNECTED_6911, SV2V_UNCONNECTED_6912, SV2V_UNCONNECTED_6913, SV2V_UNCONNECTED_6914, SV2V_UNCONNECTED_6915, SV2V_UNCONNECTED_6916, SV2V_UNCONNECTED_6917, SV2V_UNCONNECTED_6918, SV2V_UNCONNECTED_6919, SV2V_UNCONNECTED_6920, SV2V_UNCONNECTED_6921, SV2V_UNCONNECTED_6922, SV2V_UNCONNECTED_6923, SV2V_UNCONNECTED_6924, SV2V_UNCONNECTED_6925, SV2V_UNCONNECTED_6926, SV2V_UNCONNECTED_6927, SV2V_UNCONNECTED_6928, SV2V_UNCONNECTED_6929, SV2V_UNCONNECTED_6930, SV2V_UNCONNECTED_6931, SV2V_UNCONNECTED_6932, SV2V_UNCONNECTED_6933, SV2V_UNCONNECTED_6934, SV2V_UNCONNECTED_6935, SV2V_UNCONNECTED_6936, SV2V_UNCONNECTED_6937, SV2V_UNCONNECTED_6938, SV2V_UNCONNECTED_6939, SV2V_UNCONNECTED_6940, SV2V_UNCONNECTED_6941, SV2V_UNCONNECTED_6942, SV2V_UNCONNECTED_6943, SV2V_UNCONNECTED_6944, SV2V_UNCONNECTED_6945, SV2V_UNCONNECTED_6946, SV2V_UNCONNECTED_6947, SV2V_UNCONNECTED_6948, SV2V_UNCONNECTED_6949, SV2V_UNCONNECTED_6950, SV2V_UNCONNECTED_6951, SV2V_UNCONNECTED_6952, SV2V_UNCONNECTED_6953, SV2V_UNCONNECTED_6954, SV2V_UNCONNECTED_6955, SV2V_UNCONNECTED_6956, SV2V_UNCONNECTED_6957, SV2V_UNCONNECTED_6958, SV2V_UNCONNECTED_6959, SV2V_UNCONNECTED_6960, SV2V_UNCONNECTED_6961, SV2V_UNCONNECTED_6962, SV2V_UNCONNECTED_6963, SV2V_UNCONNECTED_6964, SV2V_UNCONNECTED_6965, SV2V_UNCONNECTED_6966, SV2V_UNCONNECTED_6967, SV2V_UNCONNECTED_6968, SV2V_UNCONNECTED_6969, SV2V_UNCONNECTED_6970, SV2V_UNCONNECTED_6971, SV2V_UNCONNECTED_6972, SV2V_UNCONNECTED_6973, SV2V_UNCONNECTED_6974, SV2V_UNCONNECTED_6975, SV2V_UNCONNECTED_6976, SV2V_UNCONNECTED_6977, SV2V_UNCONNECTED_6978, SV2V_UNCONNECTED_6979, SV2V_UNCONNECTED_6980, SV2V_UNCONNECTED_6981, SV2V_UNCONNECTED_6982, SV2V_UNCONNECTED_6983, SV2V_UNCONNECTED_6984, SV2V_UNCONNECTED_6985, SV2V_UNCONNECTED_6986, SV2V_UNCONNECTED_6987, SV2V_UNCONNECTED_6988, SV2V_UNCONNECTED_6989, SV2V_UNCONNECTED_6990, SV2V_UNCONNECTED_6991, SV2V_UNCONNECTED_6992, SV2V_UNCONNECTED_6993, SV2V_UNCONNECTED_6994, SV2V_UNCONNECTED_6995, SV2V_UNCONNECTED_6996, SV2V_UNCONNECTED_6997, SV2V_UNCONNECTED_6998, SV2V_UNCONNECTED_6999, SV2V_UNCONNECTED_7000, SV2V_UNCONNECTED_7001, SV2V_UNCONNECTED_7002, SV2V_UNCONNECTED_7003, SV2V_UNCONNECTED_7004, SV2V_UNCONNECTED_7005, SV2V_UNCONNECTED_7006, SV2V_UNCONNECTED_7007, SV2V_UNCONNECTED_7008, SV2V_UNCONNECTED_7009, SV2V_UNCONNECTED_7010, SV2V_UNCONNECTED_7011, SV2V_UNCONNECTED_7012, SV2V_UNCONNECTED_7013, SV2V_UNCONNECTED_7014, SV2V_UNCONNECTED_7015, SV2V_UNCONNECTED_7016, SV2V_UNCONNECTED_7017, SV2V_UNCONNECTED_7018, SV2V_UNCONNECTED_7019, SV2V_UNCONNECTED_7020, SV2V_UNCONNECTED_7021, SV2V_UNCONNECTED_7022, SV2V_UNCONNECTED_7023, SV2V_UNCONNECTED_7024, SV2V_UNCONNECTED_7025, SV2V_UNCONNECTED_7026, SV2V_UNCONNECTED_7027, SV2V_UNCONNECTED_7028, SV2V_UNCONNECTED_7029, SV2V_UNCONNECTED_7030, SV2V_UNCONNECTED_7031, SV2V_UNCONNECTED_7032, SV2V_UNCONNECTED_7033, SV2V_UNCONNECTED_7034, SV2V_UNCONNECTED_7035, SV2V_UNCONNECTED_7036, SV2V_UNCONNECTED_7037, SV2V_UNCONNECTED_7038, SV2V_UNCONNECTED_7039, SV2V_UNCONNECTED_7040, SV2V_UNCONNECTED_7041, SV2V_UNCONNECTED_7042, SV2V_UNCONNECTED_7043, SV2V_UNCONNECTED_7044, SV2V_UNCONNECTED_7045, SV2V_UNCONNECTED_7046, SV2V_UNCONNECTED_7047, SV2V_UNCONNECTED_7048, SV2V_UNCONNECTED_7049, SV2V_UNCONNECTED_7050, SV2V_UNCONNECTED_7051, SV2V_UNCONNECTED_7052, SV2V_UNCONNECTED_7053, SV2V_UNCONNECTED_7054, SV2V_UNCONNECTED_7055, SV2V_UNCONNECTED_7056, SV2V_UNCONNECTED_7057, SV2V_UNCONNECTED_7058, SV2V_UNCONNECTED_7059, SV2V_UNCONNECTED_7060, SV2V_UNCONNECTED_7061, SV2V_UNCONNECTED_7062, SV2V_UNCONNECTED_7063, SV2V_UNCONNECTED_7064, SV2V_UNCONNECTED_7065, SV2V_UNCONNECTED_7066, SV2V_UNCONNECTED_7067, SV2V_UNCONNECTED_7068, SV2V_UNCONNECTED_7069, SV2V_UNCONNECTED_7070, SV2V_UNCONNECTED_7071, SV2V_UNCONNECTED_7072, SV2V_UNCONNECTED_7073, SV2V_UNCONNECTED_7074, SV2V_UNCONNECTED_7075, SV2V_UNCONNECTED_7076, SV2V_UNCONNECTED_7077, SV2V_UNCONNECTED_7078, SV2V_UNCONNECTED_7079, SV2V_UNCONNECTED_7080, SV2V_UNCONNECTED_7081, SV2V_UNCONNECTED_7082, SV2V_UNCONNECTED_7083, SV2V_UNCONNECTED_7084, SV2V_UNCONNECTED_7085, SV2V_UNCONNECTED_7086, SV2V_UNCONNECTED_7087, SV2V_UNCONNECTED_7088, SV2V_UNCONNECTED_7089, SV2V_UNCONNECTED_7090, SV2V_UNCONNECTED_7091, SV2V_UNCONNECTED_7092, SV2V_UNCONNECTED_7093, SV2V_UNCONNECTED_7094, SV2V_UNCONNECTED_7095, SV2V_UNCONNECTED_7096, SV2V_UNCONNECTED_7097, SV2V_UNCONNECTED_7098, SV2V_UNCONNECTED_7099, SV2V_UNCONNECTED_7100, SV2V_UNCONNECTED_7101, SV2V_UNCONNECTED_7102, SV2V_UNCONNECTED_7103, SV2V_UNCONNECTED_7104, SV2V_UNCONNECTED_7105, SV2V_UNCONNECTED_7106, SV2V_UNCONNECTED_7107, SV2V_UNCONNECTED_7108, SV2V_UNCONNECTED_7109, SV2V_UNCONNECTED_7110, SV2V_UNCONNECTED_7111, SV2V_UNCONNECTED_7112, SV2V_UNCONNECTED_7113, SV2V_UNCONNECTED_7114, SV2V_UNCONNECTED_7115, SV2V_UNCONNECTED_7116, SV2V_UNCONNECTED_7117, SV2V_UNCONNECTED_7118, SV2V_UNCONNECTED_7119, SV2V_UNCONNECTED_7120, SV2V_UNCONNECTED_7121, SV2V_UNCONNECTED_7122, SV2V_UNCONNECTED_7123, SV2V_UNCONNECTED_7124, SV2V_UNCONNECTED_7125, SV2V_UNCONNECTED_7126, SV2V_UNCONNECTED_7127, SV2V_UNCONNECTED_7128, SV2V_UNCONNECTED_7129, SV2V_UNCONNECTED_7130, SV2V_UNCONNECTED_7131, SV2V_UNCONNECTED_7132, SV2V_UNCONNECTED_7133, SV2V_UNCONNECTED_7134, SV2V_UNCONNECTED_7135, SV2V_UNCONNECTED_7136, SV2V_UNCONNECTED_7137, SV2V_UNCONNECTED_7138, SV2V_UNCONNECTED_7139, SV2V_UNCONNECTED_7140, SV2V_UNCONNECTED_7141, SV2V_UNCONNECTED_7142, SV2V_UNCONNECTED_7143, SV2V_UNCONNECTED_7144, SV2V_UNCONNECTED_7145, SV2V_UNCONNECTED_7146, SV2V_UNCONNECTED_7147, SV2V_UNCONNECTED_7148, SV2V_UNCONNECTED_7149, SV2V_UNCONNECTED_7150, SV2V_UNCONNECTED_7151, SV2V_UNCONNECTED_7152, SV2V_UNCONNECTED_7153, SV2V_UNCONNECTED_7154, SV2V_UNCONNECTED_7155, SV2V_UNCONNECTED_7156, SV2V_UNCONNECTED_7157, SV2V_UNCONNECTED_7158, SV2V_UNCONNECTED_7159, SV2V_UNCONNECTED_7160, SV2V_UNCONNECTED_7161, SV2V_UNCONNECTED_7162, SV2V_UNCONNECTED_7163, SV2V_UNCONNECTED_7164, SV2V_UNCONNECTED_7165, SV2V_UNCONNECTED_7166, roundMask_E[0:0], T586, T587, T588 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> T590;
  assign N494 = ~cycleNum_B[2];
  assign N495 = N494 | cycleNum_B[3];
  assign N496 = cycleNum_B[1] | N495;
  assign N497 = N300 | N496;
  assign N498 = ~N497;
  assign N499 = N494 | cycleNum_B[3];
  assign N500 = N295 | N499;
  assign N501 = cycleNum_B[0] | N500;
  assign N502 = ~N501;
  assign N503 = N494 | cycleNum_B[3];
  assign N504 = N295 | N503;
  assign N505 = N300 | N504;
  assign N506 = ~N505;
  assign N507 = N282 | cycleNum_C[2];
  assign N508 = N309 | N507;
  assign N509 = ~N508;
  assign N510 = N494 | cycleNum_B[3];
  assign N511 = cycleNum_B[1] | N510;
  assign N512 = cycleNum_B[0] | N511;
  assign N513 = ~N512;
  assign N514 = cycleNum_E[1] | cycleNum_E[2];
  assign N515 = N286 | N514;
  assign N516 = ~N515;
  assign N517 = T137[0] | T137[1];
  assign N518 = specialCodeB_PA[0] | N517;
  assign N519 = ~N518;
  assign N520 = T139[0] | T139[1];
  assign N521 = specialCodeA_PA[0] | N520;
  assign N522 = ~N521;
  assign N523 = T139[0] & T139[1];
  assign N524 = T137[0] & T137[1];
  assign N525 = T114[0] | T114[1];
  assign N526 = specialCodeB_PB[0] | N525;
  assign N527 = ~N526;
  assign N528 = T116[0] | T116[1];
  assign N529 = specialCodeA_PB[0] | N528;
  assign N530 = ~N529;
  assign N531 = T51[0] | T51[1];
  assign N532 = specialCodeB_PC[0] | N531;
  assign N533 = ~N532;
  assign N534 = T53[0] | T53[1];
  assign N535 = specialCodeA_PC[0] | N534;
  assign N536 = ~N535;
  assign N537 = T116[0] & T116[1];
  assign N538 = T114[0] & T114[1];
  assign N539 = T53[0] & T53[1];
  assign N540 = T51[0] & T51[1];
  assign { T198_13, T198[11:11] } = 1'b0 - io_b[63];
  assign T29 = cycleNum_E - 1'b1;
  assign T72 = cycleNum_C - 1'b1;
  assign T77 = cycleNum_B - 1'b1;
  assign T82 = cycleNum_A - 1'b1;
  assign T284 = T285 + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign T592 = T593 + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { T598, expP2_PC[0:0] } = { T593, exp_PC[0:0] } + { 1'b1, 1'b0 };
  assign T302 = { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } + { T256, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign T197 = io_a[63:52] + { T198_13, T198_13, T198 };
  assign T711 = T598 + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { T339[5:5], T339_0 } = 1'b0 - N349;
  assign sigAdjT_E = T727 + T944[0];
  assign { sigY1_E_53, SV2V_UNCONNECTED_7167, sigY1_E } = T728 + 1'b1;
  assign { T305[7:7], T305_0 } = 1'b0 - T305[20];
  assign T916 = mulAdd9A_A * mulAdd9B_A;
  assign T461 = mulAdd9C_A + 1'b1;
  assign { loMulAdd9Out_A[18:18], T251[8:0], mulAdd9Out_A } = T916 + T253;
  assign { T817[51:51], T817_0 } = 1'b0 - T946[0];
  assign T885 = (N0)? T2 : 
                (N1)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = cyc_E3_sqrt;
  assign N1 = N119;
  assign T9 = (N2)? T10 : 
              (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = T13;
  assign N3 = N120;
  assign T17 = (N4)? sqrtOp_PB : 
               (N5)? io_sqrtOp : 1'b0;
  assign N4 = valid_PB;
  assign N5 = N121;
  assign T19 = (N6)? sqrtOp_PA : 
               (N7)? io_sqrtOp : 1'b0;
  assign N6 = valid_PA;
  assign N7 = N122;
  assign valid_leaving_PB = (N8)? N509 : 
                            (N9)? ready_PC : 1'b0;
  assign N8 = normalCase_PB;
  assign N9 = N123;
  assign T28 = (N10)? { 1'b1, 1'b0, 1'b0 } : 
               (N11)? T29 : 1'b0;
  assign N10 = N312;
  assign N11 = N311;
  assign normalCase_PC = (N12)? T54 : 
                         (N13)? T33 : 1'b0;
  assign N12 = sqrtOp_PC;
  assign N13 = N124;
  assign T36 = (N4)? { T114, specialCodeB_PB[0:0] } : 
               (N5)? io_b[63:61] : 1'b0;
  assign T38 = (N6)? { T137, specialCodeB_PA[0:0] } : 
               (N7)? io_b[63:61] : 1'b0;
  assign T43 = (N4)? { T116, specialCodeA_PB[0:0] } : 
               (N5)? io_a[63:61] : 1'b0;
  assign T45 = (N6)? { T139, specialCodeA_PA[0:0] } : 
               (N7)? io_a[63:61] : 1'b0;
  assign T57 = (N4)? sign_PB : 
               (N5)? sign_S : 1'b0;
  assign sign_S = (N14)? io_b[64] : 
                  (N15)? T58 : 1'b0;
  assign N14 = io_sqrtOp;
  assign N15 = N131;
  assign T60 = (N6)? sign_PA : 
               (N7)? sign_S : 1'b0;
  assign T71 = (N16)? { 1'b1, T73 } : 
               (N17)? T72 : 1'b0;
  assign N16 = N489;
  assign N17 = N488;
  assign T76 = (N18)? { T78, 1'b1, 1'b0 } : 
               (N19)? T77 : 1'b0;
  assign N18 = T475[51];
  assign N19 = N315;
  assign T81 = (N20)? T82 : 
               (N21)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = T83;
  assign N21 = N127;
  assign normalCase_PB = (N22)? T117 : 
                         (N23)? T108 : 1'b0;
  assign N22 = sqrtOp_PB;
  assign N23 = N125;
  assign valid_leaving_PA = (N24)? valid_normalCase_leaving_PA : 
                            (N25)? ready_PB : 1'b0;
  assign N24 = normalCase_PA;
  assign N25 = N128;
  assign normalCase_PA = (N26)? T140 : 
                         (N27)? T131 : 1'b0;
  assign N26 = sqrtOp_PA;
  assign N27 = N126;
  assign normalCase_S = (N14)? normalCase_S_sqrt : 
                        (N15)? normalCase_S_div : 1'b0;
  assign T162 = (N28)? T163 : 
                (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = T165;
  assign N29 = N129;
  assign T169 = (N30)? { T170[0:0], 1'b0 } : 
                (N31)? T170 : 1'b0;
  assign N30 = exp_PC[0];
  assign N31 = N130;
  assign T180 = (N4)? fractB_51_PB : 
                (N5)? io_b[51] : 1'b0;
  assign T183 = (N6)? sigB_PA_51 : 
                (N7)? io_b[51] : 1'b0;
  assign T196 = (N14)? { 1'b0, 1'b0, io_b[63:52] } : 
                (N15)? T197 : 1'b0;
  assign T897[53] = (N32)? T206[53] : 
                    (N33)? 1'b0 : 1'b0;
  assign N32 = T212;
  assign N33 = N132;
  assign T217 = (N34)? T218 : 
                (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = T225;
  assign N35 = N133;
  assign T898 = (N36)? T230 : 
                (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = N308;
  assign N37 = N307;
  assign T233 = (N16)? T230 : 
                (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T900 = (N38)? { sqrSigma1_C, T241, sqrSigma1_C_0 } : 
                (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = N476;
  assign N39 = N475;
  assign T901 = (N36)? T241 : 
                (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T902 = (N40)? T244 : 
                (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N513;
  assign N41 = N512;
  assign T247 = (N42)? T248 : 
                (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = cyc_B6_sqrt;
  assign N43 = N134;
  assign ER1_A1_sqrt[15:0] = (N44)? { T903, 1'b0 } : 
                             (N45)? { 1'b1, T903 } : 1'b0;
  assign N44 = ER1_A1_sqrt[16];
  assign N45 = N135;
  assign T903 = (N26)? T251[15:1] : 
                (N27)? T251[14:0] : 1'b0;
  assign T904 = (N46)? T256 : 
                (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = cyc_A1_div;
  assign N47 = N136;
  assign zFractR0_A4_div = (N48)? T260 : 
                           (N49)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = T262;
  assign N49 = N137;
  assign zFractR0_A6_sqrt = (N50)? T265 : 
                            (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = T267;
  assign N51 = N138;
  assign T272 = (N52)? T256 : 
                (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = cyc_A1_sqrt;
  assign N53 = N139;
  assign T275 = (N54)? partNegSigma0_A : 
                (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = T281;
  assign N55 = N140;
  assign T277 = (N56)? { T251[11:0], mulAdd9Out_A } : 
                (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T251 } : 1'b0;
  assign N56 = N327;
  assign N57 = N326;
  assign T283 = (N58)? T284 : 
                (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = T287;
  assign N59 = N141;
  assign { T292, sqrR0_A5_sqrt } = (N60)? { T251[9:0], mulAdd9Out_A } : 
                                   (N45)? { T251[10:0], mulAdd9Out_A[8:1] } : 1'b0;
  assign N60 = exp_PA[0];
  assign T911 = (N61)? T302 : 
                (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N61 = N324;
  assign N62 = N323;
  assign T388 = (N63)? nextMulAdd9B_A : 
                (N64)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N63 = T407;
  assign N64 = N142;
  assign T391[7:0] = (N65)? T256[23:16] : 
                     (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N65 = T391[8];
  assign N66 = N319;
  assign T395 = (N56)? T908[8:0] : 
                (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T399 = (N61)? sqrR0_A5_sqrt : 
                (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T402 = (N67)? io_b[50:42] : 
                (N68)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = cyc_A7_sqrt;
  assign N68 = N143;
  assign T424 = (N69)? T918 : 
                (N70)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N69 = T450;
  assign N70 = N144;
  assign T917 = (N71)? T426 : 
                (N72)? T918 : 1'b0;
  assign N71 = T445;
  assign N72 = N145;
  assign T919 = (N73)? T428 : 
                (N74)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N73 = T430;
  assign N74 = N146;
  assign T920[7:0] = (N75)? { sigB_PA_51, sigB_PA_50, sigB_PA_49, sigB_PA_48, sigB_PA_47, T285[20:18] } : 
                     (N76)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N75 = T920[8];
  assign N76 = N147;
  assign { zFractB_A4_div, T921 } = (N77)? io_b[48:35] : 
                                    (N78)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N77 = T305[20];
  assign N78 = N148;
  assign T922 = (N56)? T285[17:9] : 
                (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T442 = (N67)? T443 : 
                (N68)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T251[15:9] = (N79)? T461 : 
                      (N80)? mulAdd9C_A : 1'b0;
  assign N79 = loMulAdd9Out_A[18];
  assign N80 = N149;
  assign T926 = (N81)? T472 : 
                (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N81 = N506;
  assign N82 = N505;
  assign T475[50:36] = (N18)? T903 : 
                       (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign zComplSigT_C1_sqrt = (N83)? T485 : 
                              (N84)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N83 = cyc_C1_sqrt;
  assign N84 = N150;
  assign T488[51:0] = (N85)? { sigB_PC, T170[0:0] } : 
                      (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N85 = T488[52];
  assign N86 = N151;
  assign T928 = (N87)? T491 : 
                (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N87 = cyc_C4_sqrt;
  assign N88 = N152;
  assign T929 = (N89)? T218[104:72] : 
                (N90)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N89 = cyc_C4_div;
  assign N90 = N153;
  assign T930 = (N91)? io_mulAddResult_3[104:59] : 
                (N92)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N91 = T502;
  assign N92 = N154;
  assign T506[51:0] = (N93)? sigA_PA : 
                      (N94)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N93 = T506[52];
  assign N94 = N155;
  assign T514[51:0] = (N95)? { sigB_PA_51, sigB_PA_50, sigB_PA_49, sigB_PA_48, sigB_PA_47, T285, sigB_PA } : 
                      (N96)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N95 = T514[52];
  assign N96 = N156;
  assign T516 = (N52)? ER1_A1_sqrt : 
                (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T933 = (N12)? T592 : 
                (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T595 = (N97)? expP1_PC : 
                (N98)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N97 = T601;
  assign N98 = N157;
  assign expP1_PC[13:1] = (N30)? T598 : 
                          (N99)? T593 : 1'b0;
  assign N99 = expP1_PC[0];
  assign T604 = (N100)? { T593, exp_PC[0:0] } : 
                (N101)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N100 = T605;
  assign N101 = N158;
  assign trueLtX_E1 = (N12)? T696 : 
                      (N13)? isNegRemT_E : 1'b0;
  assign T693 = (N12)? io_mulAddResult_3[55] : 
                (N13)? io_mulAddResult_3[53] : 1'b0;
  assign T943 = (N102)? T711 : 
                (N103)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N102 = T713;
  assign N103 = N159;
  assign { roundEvenMask_E1_53, roundEvenMask_E1 } = (N104)? { T701[52:52], T701[50:0], incrPosMask_E[0:0] } : 
                                                     (N105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N104 = T716;
  assign N105 = N160;
  assign T720 = (N4)? roundingMode_PB : 
                (N5)? io_roundingMode : 1'b0;
  assign T722 = (N6)? roundingMode_PA : 
                (N7)? io_roundingMode : 1'b0;
  assign { T724_53, T724 } = (N106)? { sigY1_E_53, sigY1_E } : 
                             (N107)? { sigY0_E_53, sigY0_E } : 1'b0;
  assign N106 = T730;
  assign N107 = N161;
  assign T944[0] = (N108)? N469 : 
                   (N109)? N470 : 1'b0;
  assign N108 = sign_PC;
  assign N109 = N162;
  assign T760 = (N110)? { T598, expP2_PC[0:0] } : 
                (N111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N110 = T761;
  assign N111 = N163;
  assign T767 = (N112)? expP1_PC : 
                (N113)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N112 = T768;
  assign N113 = N164;
  assign T772 = (N114)? { sExpX_E[13:13], posExpX_E } : 
                (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N114 = T773;
  assign N115 = N165;
  assign notSigNaN_invalid_PC = (N12)? T793 : 
                                (N13)? T786 : 1'b0;
  assign T803 = (N4)? fractA_51_PB : 
                (N5)? io_a[51] : 1'b0;
  assign T806 = (N6)? sigA_PA[51] : 
                (N7)? io_a[51] : 1'b0;
  assign T819 = (N116)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N117)? sigY_E1 : 1'b0;
  assign N116 = T820;
  assign N117 = N166;
  assign notSpecial_isZeroOut_E1 = (N12)? N533 : 
                                   (N13)? T822 : 1'b0;
  assign notNaN_isInfOut_E1 = (N12)? isInfB_PC : 
                              (N13)? T829 : 1'b0;
  assign T849 = (N12)? T850 : 
                (N13)? sign_PC : 1'b0;
  assign N169 = (N118)? 1'b1 : 
                (N205)? 1'b1 : 
                (N168)? 1'b0 : 1'b0;
  assign N118 = reset;
  assign { N172, N171, N170 } = (N118)? { 1'b0, 1'b0, 1'b0 } : 
                                (N205)? T28 : 1'b0;
  assign N175 = (N118)? 1'b1 : 
                (N206)? 1'b1 : 
                (N174)? 1'b0 : 1'b0;
  assign N176 = (N118)? 1'b0 : 
                (N206)? entering_PC : 1'b0;
  assign N179 = (N118)? 1'b1 : 
                (N207)? 1'b1 : 
                (N178)? 1'b0 : 1'b0;
  assign { N182, N181, N180 } = (N118)? { 1'b0, 1'b0, 1'b0 } : 
                                (N207)? T71 : 1'b0;
  assign N185 = (N118)? 1'b1 : 
                (N208)? 1'b1 : 
                (N184)? 1'b0 : 1'b0;
  assign { N189, N188, N187, N186 } = (N118)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N208)? T76 : 1'b0;
  assign N192 = (N118)? 1'b1 : 
                (N209)? 1'b1 : 
                (N191)? 1'b0 : 1'b0;
  assign { N195, N194, N193 } = (N118)? { 1'b0, 1'b0, 1'b0 } : 
                                (N209)? T80 : 1'b0;
  assign N198 = (N118)? 1'b1 : 
                (N210)? 1'b1 : 
                (N197)? 1'b0 : 1'b0;
  assign N199 = (N118)? 1'b0 : 
                (N210)? entering_PA : 1'b0;
  assign N202 = (N118)? 1'b1 : 
                (N211)? 1'b1 : 
                (N201)? 1'b0 : 1'b0;
  assign N203 = (N118)? 1'b0 : 
                (N211)? entering_PB : 1'b0;
  assign io_mulAddC_2[104] = T204[104] | 1'b0;
  assign io_mulAddC_2[103] = T204[103] | 1'b0;
  assign io_mulAddC_2[102] = T204[102] | 1'b0;
  assign io_mulAddC_2[101] = T204[101] | 1'b0;
  assign io_mulAddC_2[100] = T204[100] | 1'b0;
  assign io_mulAddC_2[99] = T204[99] | 1'b0;
  assign io_mulAddC_2[98] = T204[98] | 1'b0;
  assign io_mulAddC_2[97] = T204[97] | 1'b0;
  assign io_mulAddC_2[96] = T204[96] | 1'b0;
  assign io_mulAddC_2[95] = T204[95] | 1'b0;
  assign io_mulAddC_2[94] = T204[94] | 1'b0;
  assign io_mulAddC_2[93] = T204[93] | 1'b0;
  assign io_mulAddC_2[92] = T204[92] | 1'b0;
  assign io_mulAddC_2[91] = T204[91] | 1'b0;
  assign io_mulAddC_2[90] = T204[90] | 1'b0;
  assign io_mulAddC_2[89] = T204[89] | 1'b0;
  assign io_mulAddC_2[88] = T204[88] | 1'b0;
  assign io_mulAddC_2[87] = T204[87] | 1'b0;
  assign io_mulAddC_2[86] = T204[86] | 1'b0;
  assign io_mulAddC_2[85] = T204[85] | 1'b0;
  assign io_mulAddC_2[84] = T204[84] | 1'b0;
  assign io_mulAddC_2[83] = T204[83] | 1'b0;
  assign io_mulAddC_2[82] = T204[82] | 1'b0;
  assign io_mulAddC_2[81] = T204[81] | 1'b0;
  assign io_mulAddC_2[80] = T204[80] | 1'b0;
  assign io_mulAddC_2[79] = T204[79] | 1'b0;
  assign io_mulAddC_2[78] = T204[78] | 1'b0;
  assign io_mulAddC_2[77] = T204[77] | 1'b0;
  assign io_mulAddC_2[76] = T204[76] | 1'b0;
  assign io_mulAddC_2[75] = T204[75] | 1'b0;
  assign io_mulAddC_2[74] = T204[74] | 1'b0;
  assign io_mulAddC_2[73] = T204[73] | 1'b0;
  assign io_mulAddC_2[72] = T204[72] | 1'b0;
  assign io_mulAddC_2[71] = T204[71] | 1'b0;
  assign io_mulAddC_2[70] = T204[70] | 1'b0;
  assign io_mulAddC_2[69] = T204[69] | 1'b0;
  assign io_mulAddC_2[68] = T204[68] | 1'b0;
  assign io_mulAddC_2[67] = T204[67] | 1'b0;
  assign io_mulAddC_2[66] = T204[66] | 1'b0;
  assign io_mulAddC_2[65] = T204[65] | 1'b0;
  assign io_mulAddC_2[64] = T204[64] | 1'b0;
  assign io_mulAddC_2[63] = T204[63] | 1'b0;
  assign io_mulAddC_2[62] = T204[62] | 1'b0;
  assign io_mulAddC_2[61] = T204[61] | 1'b0;
  assign io_mulAddC_2[60] = T204[60] | 1'b0;
  assign io_mulAddC_2[59] = T204[59] | 1'b0;
  assign io_mulAddC_2[58] = T204[58] | 1'b0;
  assign io_mulAddC_2[57] = T204[57] | 1'b0;
  assign io_mulAddC_2[56] = T204[56] | 1'b0;
  assign io_mulAddC_2[55] = T204[55] | T885[55];
  assign io_mulAddC_2[54] = T204[54] | T885[54];
  assign io_mulAddC_2[53] = T204[53] | 1'b0;
  assign io_mulAddC_2[52] = T204[52] | 1'b0;
  assign io_mulAddC_2[51] = T204[51] | 1'b0;
  assign io_mulAddC_2[50] = T204[50] | 1'b0;
  assign io_mulAddC_2[49] = T204[49] | 1'b0;
  assign io_mulAddC_2[48] = T204[48] | 1'b0;
  assign io_mulAddC_2[47] = T204[47] | 1'b0;
  assign io_mulAddC_2[46] = T204[46] | 1'b0;
  assign io_mulAddC_2[45] = T204[45] | 1'b0;
  assign io_mulAddC_2[44] = T204[44] | 1'b0;
  assign io_mulAddC_2[43] = T204[43] | 1'b0;
  assign io_mulAddC_2[42] = T204[42] | 1'b0;
  assign io_mulAddC_2[41] = T204[41] | 1'b0;
  assign io_mulAddC_2[40] = T204[40] | 1'b0;
  assign io_mulAddC_2[39] = T204[39] | 1'b0;
  assign io_mulAddC_2[38] = T204[38] | 1'b0;
  assign io_mulAddC_2[37] = T204[37] | 1'b0;
  assign io_mulAddC_2[36] = T204[36] | 1'b0;
  assign io_mulAddC_2[35] = T204[35] | 1'b0;
  assign io_mulAddC_2[34] = T204[34] | 1'b0;
  assign io_mulAddC_2[33] = T204[33] | 1'b0;
  assign io_mulAddC_2[32] = T204[32] | 1'b0;
  assign io_mulAddC_2[31] = T204[31] | 1'b0;
  assign io_mulAddC_2[30] = T204[30] | 1'b0;
  assign io_mulAddC_2[29] = T204[29] | 1'b0;
  assign io_mulAddC_2[28] = T204[28] | 1'b0;
  assign io_mulAddC_2[27] = T204[27] | 1'b0;
  assign io_mulAddC_2[26] = T204[26] | 1'b0;
  assign io_mulAddC_2[25] = T204[25] | 1'b0;
  assign io_mulAddC_2[24] = T204[24] | 1'b0;
  assign io_mulAddC_2[23] = T204[23] | 1'b0;
  assign io_mulAddC_2[22] = T204[22] | 1'b0;
  assign io_mulAddC_2[21] = T204[21] | 1'b0;
  assign io_mulAddC_2[20] = T204[20] | 1'b0;
  assign io_mulAddC_2[19] = T204[19] | 1'b0;
  assign io_mulAddC_2[18] = T204[18] | 1'b0;
  assign io_mulAddC_2[17] = T204[17] | 1'b0;
  assign io_mulAddC_2[16] = T204[16] | 1'b0;
  assign io_mulAddC_2[15] = T204[15] | 1'b0;
  assign io_mulAddC_2[14] = T204[14] | 1'b0;
  assign io_mulAddC_2[13] = T204[13] | 1'b0;
  assign io_mulAddC_2[12] = T204[12] | 1'b0;
  assign io_mulAddC_2[11] = T204[11] | 1'b0;
  assign io_mulAddC_2[10] = T204[10] | 1'b0;
  assign io_mulAddC_2[9] = T204[9] | 1'b0;
  assign io_mulAddC_2[8] = T204[8] | 1'b0;
  assign io_mulAddC_2[7] = T204[7] | 1'b0;
  assign io_mulAddC_2[6] = T204[6] | 1'b0;
  assign io_mulAddC_2[5] = T204[5] | 1'b0;
  assign io_mulAddC_2[4] = T204[4] | 1'b0;
  assign io_mulAddC_2[3] = T204[3] | 1'b0;
  assign io_mulAddC_2[2] = T204[2] | 1'b0;
  assign io_mulAddC_2[1] = T204[1] | 1'b0;
  assign io_mulAddC_2[0] = T204[0] | 1'b0;
  assign N119 = ~cyc_E3_sqrt;
  assign T2[55] = T169[1] ^ T4[1];
  assign T2[54] = T169[0] ^ 1'b0;
  assign T4[1] = ~extraT_E;
  assign sigT_C1[53] = ~zComplSigT_C1[53];
  assign sigT_C1[52] = ~zComplSigT_C1[52];
  assign sigT_C1[51] = ~zComplSigT_C1[51];
  assign sigT_C1[50] = ~zComplSigT_C1[50];
  assign sigT_C1[49] = ~zComplSigT_C1[49];
  assign sigT_C1[48] = ~zComplSigT_C1[48];
  assign sigT_C1[47] = ~zComplSigT_C1[47];
  assign sigT_C1[46] = ~zComplSigT_C1[46];
  assign sigT_C1[45] = ~zComplSigT_C1[45];
  assign sigT_C1[44] = ~zComplSigT_C1[44];
  assign sigT_C1[43] = ~zComplSigT_C1[43];
  assign sigT_C1[42] = ~zComplSigT_C1[42];
  assign sigT_C1[41] = ~zComplSigT_C1[41];
  assign sigT_C1[40] = ~zComplSigT_C1[40];
  assign sigT_C1[39] = ~zComplSigT_C1[39];
  assign sigT_C1[38] = ~zComplSigT_C1[38];
  assign sigT_C1[37] = ~zComplSigT_C1[37];
  assign sigT_C1[36] = ~zComplSigT_C1[36];
  assign sigT_C1[35] = ~zComplSigT_C1[35];
  assign sigT_C1[34] = ~zComplSigT_C1[34];
  assign sigT_C1[33] = ~zComplSigT_C1[33];
  assign sigT_C1[32] = ~zComplSigT_C1[32];
  assign sigT_C1[31] = ~zComplSigT_C1[31];
  assign sigT_C1[30] = ~zComplSigT_C1[30];
  assign sigT_C1[29] = ~zComplSigT_C1[29];
  assign sigT_C1[28] = ~zComplSigT_C1[28];
  assign sigT_C1[27] = ~zComplSigT_C1[27];
  assign sigT_C1[26] = ~zComplSigT_C1[26];
  assign sigT_C1[25] = ~zComplSigT_C1[25];
  assign sigT_C1[24] = ~zComplSigT_C1[24];
  assign sigT_C1[23] = ~zComplSigT_C1[23];
  assign sigT_C1[22] = ~zComplSigT_C1[22];
  assign sigT_C1[21] = ~zComplSigT_C1[21];
  assign sigT_C1[20] = ~zComplSigT_C1[20];
  assign sigT_C1[19] = ~zComplSigT_C1[19];
  assign sigT_C1[18] = ~zComplSigT_C1[18];
  assign sigT_C1[17] = ~zComplSigT_C1[17];
  assign sigT_C1[16] = ~zComplSigT_C1[16];
  assign sigT_C1[15] = ~zComplSigT_C1[15];
  assign sigT_C1[14] = ~zComplSigT_C1[14];
  assign sigT_C1[13] = ~zComplSigT_C1[13];
  assign sigT_C1[12] = ~zComplSigT_C1[12];
  assign sigT_C1[11] = ~zComplSigT_C1[11];
  assign sigT_C1[10] = ~zComplSigT_C1[10];
  assign sigT_C1[9] = ~zComplSigT_C1[9];
  assign sigT_C1[8] = ~zComplSigT_C1[8];
  assign sigT_C1[7] = ~zComplSigT_C1[7];
  assign sigT_C1[6] = ~zComplSigT_C1[6];
  assign sigT_C1[5] = ~zComplSigT_C1[5];
  assign sigT_C1[4] = ~zComplSigT_C1[4];
  assign sigT_C1[3] = ~zComplSigT_C1[3];
  assign sigT_C1[2] = ~zComplSigT_C1[2];
  assign sigT_C1[1] = ~zComplSigT_C1[1];
  assign sigT_C1[0] = ~zComplSigT_C1[0];
  assign zComplSigT_C1[53] = T162[53] | 1'b0;
  assign zComplSigT_C1[52] = T162[52] | T9[52];
  assign zComplSigT_C1[51] = T162[51] | T9[51];
  assign zComplSigT_C1[50] = T162[50] | T9[50];
  assign zComplSigT_C1[49] = T162[49] | T9[49];
  assign zComplSigT_C1[48] = T162[48] | T9[48];
  assign zComplSigT_C1[47] = T162[47] | T9[47];
  assign zComplSigT_C1[46] = T162[46] | T9[46];
  assign zComplSigT_C1[45] = T162[45] | T9[45];
  assign zComplSigT_C1[44] = T162[44] | T9[44];
  assign zComplSigT_C1[43] = T162[43] | T9[43];
  assign zComplSigT_C1[42] = T162[42] | T9[42];
  assign zComplSigT_C1[41] = T162[41] | T9[41];
  assign zComplSigT_C1[40] = T162[40] | T9[40];
  assign zComplSigT_C1[39] = T162[39] | T9[39];
  assign zComplSigT_C1[38] = T162[38] | T9[38];
  assign zComplSigT_C1[37] = T162[37] | T9[37];
  assign zComplSigT_C1[36] = T162[36] | T9[36];
  assign zComplSigT_C1[35] = T162[35] | T9[35];
  assign zComplSigT_C1[34] = T162[34] | T9[34];
  assign zComplSigT_C1[33] = T162[33] | T9[33];
  assign zComplSigT_C1[32] = T162[32] | T9[32];
  assign zComplSigT_C1[31] = T162[31] | T9[31];
  assign zComplSigT_C1[30] = T162[30] | T9[30];
  assign zComplSigT_C1[29] = T162[29] | T9[29];
  assign zComplSigT_C1[28] = T162[28] | T9[28];
  assign zComplSigT_C1[27] = T162[27] | T9[27];
  assign zComplSigT_C1[26] = T162[26] | T9[26];
  assign zComplSigT_C1[25] = T162[25] | T9[25];
  assign zComplSigT_C1[24] = T162[24] | T9[24];
  assign zComplSigT_C1[23] = T162[23] | T9[23];
  assign zComplSigT_C1[22] = T162[22] | T9[22];
  assign zComplSigT_C1[21] = T162[21] | T9[21];
  assign zComplSigT_C1[20] = T162[20] | T9[20];
  assign zComplSigT_C1[19] = T162[19] | T9[19];
  assign zComplSigT_C1[18] = T162[18] | T9[18];
  assign zComplSigT_C1[17] = T162[17] | T9[17];
  assign zComplSigT_C1[16] = T162[16] | T9[16];
  assign zComplSigT_C1[15] = T162[15] | T9[15];
  assign zComplSigT_C1[14] = T162[14] | T9[14];
  assign zComplSigT_C1[13] = T162[13] | T9[13];
  assign zComplSigT_C1[12] = T162[12] | T9[12];
  assign zComplSigT_C1[11] = T162[11] | T9[11];
  assign zComplSigT_C1[10] = T162[10] | T9[10];
  assign zComplSigT_C1[9] = T162[9] | T9[9];
  assign zComplSigT_C1[8] = T162[8] | T9[8];
  assign zComplSigT_C1[7] = T162[7] | T9[7];
  assign zComplSigT_C1[6] = T162[6] | T9[6];
  assign zComplSigT_C1[5] = T162[5] | T9[5];
  assign zComplSigT_C1[4] = T162[4] | T9[4];
  assign zComplSigT_C1[3] = T162[3] | T9[3];
  assign zComplSigT_C1[2] = T162[2] | T9[2];
  assign zComplSigT_C1[1] = T162[1] | T9[1];
  assign zComplSigT_C1[0] = T162[0] | T9[0];
  assign N120 = ~T13;
  assign T10[52] = ~io_mulAddResult_3[102];
  assign T10[51] = ~io_mulAddResult_3[101];
  assign T10[50] = ~io_mulAddResult_3[100];
  assign T10[49] = ~io_mulAddResult_3[99];
  assign T10[48] = ~io_mulAddResult_3[98];
  assign T10[47] = ~io_mulAddResult_3[97];
  assign T10[46] = ~io_mulAddResult_3[96];
  assign T10[45] = ~io_mulAddResult_3[95];
  assign T10[44] = ~io_mulAddResult_3[94];
  assign T10[43] = ~io_mulAddResult_3[93];
  assign T10[42] = ~io_mulAddResult_3[92];
  assign T10[41] = ~io_mulAddResult_3[91];
  assign T10[40] = ~io_mulAddResult_3[90];
  assign T10[39] = ~io_mulAddResult_3[89];
  assign T10[38] = ~io_mulAddResult_3[88];
  assign T10[37] = ~io_mulAddResult_3[87];
  assign T10[36] = ~io_mulAddResult_3[86];
  assign T10[35] = ~io_mulAddResult_3[85];
  assign T10[34] = ~io_mulAddResult_3[84];
  assign T10[33] = ~io_mulAddResult_3[83];
  assign T10[32] = ~io_mulAddResult_3[82];
  assign T10[31] = ~io_mulAddResult_3[81];
  assign T10[30] = ~io_mulAddResult_3[80];
  assign T10[29] = ~io_mulAddResult_3[79];
  assign T10[28] = ~io_mulAddResult_3[78];
  assign T10[27] = ~io_mulAddResult_3[77];
  assign T10[26] = ~io_mulAddResult_3[76];
  assign T10[25] = ~io_mulAddResult_3[75];
  assign T10[24] = ~io_mulAddResult_3[74];
  assign T10[23] = ~io_mulAddResult_3[73];
  assign T10[22] = ~io_mulAddResult_3[72];
  assign T10[21] = ~io_mulAddResult_3[71];
  assign T10[20] = ~io_mulAddResult_3[70];
  assign T10[19] = ~io_mulAddResult_3[69];
  assign T10[18] = ~io_mulAddResult_3[68];
  assign T10[17] = ~io_mulAddResult_3[67];
  assign T10[16] = ~io_mulAddResult_3[66];
  assign T10[15] = ~io_mulAddResult_3[65];
  assign T10[14] = ~io_mulAddResult_3[64];
  assign T10[13] = ~io_mulAddResult_3[63];
  assign T10[12] = ~io_mulAddResult_3[62];
  assign T10[11] = ~io_mulAddResult_3[61];
  assign T10[10] = ~io_mulAddResult_3[60];
  assign T10[9] = ~io_mulAddResult_3[59];
  assign T10[8] = ~io_mulAddResult_3[58];
  assign T10[7] = ~io_mulAddResult_3[57];
  assign T10[6] = ~io_mulAddResult_3[56];
  assign T10[5] = ~io_mulAddResult_3[55];
  assign T10[4] = ~io_mulAddResult_3[54];
  assign T10[3] = ~io_mulAddResult_3[53];
  assign T10[2] = ~io_mulAddResult_3[52];
  assign T10[1] = ~io_mulAddResult_3[51];
  assign T10[0] = ~io_mulAddResult_3[50];
  assign T13 = cyc_C1_div & E_C1_div;
  assign E_C1_div = ~io_mulAddResult_3[104];
  assign cyc_C1_div = N312 & T15;
  assign T15 = ~sqrtOp_PC;
  assign N121 = ~valid_PB;
  assign N122 = ~valid_PA;
  assign entering_PA = entering_PA_normalCase | T21;
  assign T21 = cyc_S & T22;
  assign T22 = valid_PA | T23;
  assign T23 = ~ready_PB;
  assign ready_PB = T122 | valid_leaving_PB;
  assign N123 = ~normalCase_PB;
  assign ready_PC = T65 | valid_leaving_PC;
  assign valid_leaving_PC = T32 | N516;
  assign T30 = N312 | N274;
  assign T32 = ~normalCase_PC;
  assign N124 = ~sqrtOp_PC;
  assign T33 = T40 & T34;
  assign T34 = ~N533;
  assign T40 = T49 & T41;
  assign T41 = ~N536;
  assign T47 = entering_PA & T48;
  assign T48 = ~io_sqrtOp;
  assign T49 = T52 & T50;
  assign T50 = ~N540;
  assign T52 = ~N539;
  assign T54 = T62 & T55;
  assign T55 = ~sign_PC;
  assign T58 = io_a[64] ^ io_b[64];
  assign T62 = T64 & T63;
  assign T63 = ~N533;
  assign T64 = ~N540;
  assign T65 = ~valid_PC;
  assign T67 = entering_PC | leaving_PC;
  assign leaving_PC = valid_PC & valid_leaving_PC;
  assign N125 = ~sqrtOp_PB;
  assign T73[1] = sqrtOp_PB;
  assign T73[0] = N125;
  assign T475[51] = N316;
  assign N126 = ~sqrtOp_PA;
  assign T78[3] = sqrtOp_PA;
  assign T78[2] = N126;
  assign T80[2] = T84[2] | T81[2];
  assign T80[1] = T84[1] | T81[1];
  assign T80[0] = T84[0] | T81[0];
  assign N127 = ~T83;
  assign T83 = ~entering_PA_normalCase;
  assign T84[2] = 1'b0 | T85[2];
  assign T84[1] = T891[1] | T85[2];
  assign T84[0] = T891[1] | 1'b0;
  assign T85[2] = cyc_A7_sqrt;
  assign cyc_A7_sqrt = cyc_S_sqrt & normalCase_S_sqrt;
  assign normalCase_S_sqrt = T87 & T86;
  assign T86 = ~io_b[64];
  assign T87 = T89 & T88;
  assign T88 = ~N466;
  assign T89 = ~N478;
  assign cyc_S_sqrt = T91 & io_sqrtOp;
  assign T91 = io_inReady_sqrt & io_inValid;
  assign T891[1] = T305[20];
  assign T305[20] = cyc_S_div & normalCase_S_div;
  assign normalCase_S_div = T94 & T93;
  assign T93 = ~N466;
  assign T94 = T96 & T95;
  assign T95 = ~N473;
  assign T96 = T98 & T97;
  assign T97 = ~N478;
  assign T98 = ~N477;
  assign cyc_S_div = T101 & T100;
  assign T100 = ~io_sqrtOp;
  assign T101 = io_inReady_div & io_inValid;
  assign T102 = entering_PA_normalCase | N281;
  assign T104 = N316 | N279;
  assign T106 = N489 | N276;
  assign T108 = T110 & T109;
  assign T109 = ~N527;
  assign T110 = T112 & T111;
  assign T111 = ~N530;
  assign T112 = T115 & T113;
  assign T113 = ~N538;
  assign T115 = ~N537;
  assign T117 = T119 & T118;
  assign T118 = ~sign_PB;
  assign T119 = T121 & T120;
  assign T120 = ~N527;
  assign T121 = ~N538;
  assign T122 = ~valid_PB;
  assign cyc_S = cyc_S_div | cyc_S_sqrt;
  assign entering_PA_normalCase = T305[20] | cyc_A7_sqrt;
  assign T124 = entering_PA | leaving_PA;
  assign leaving_PA = valid_PA & valid_leaving_PA;
  assign N128 = ~normalCase_PA;
  assign valid_normalCase_leaving_PA = cyc_B4_div | N506;
  assign cyc_B4_div = T129 & T128;
  assign T128 = ~sqrtOp_PA;
  assign T129 = N513 & valid_PA;
  assign T131 = T133 & T132;
  assign T132 = ~N519;
  assign T133 = T135 & T134;
  assign T134 = ~N522;
  assign T135 = T138 & T136;
  assign T136 = ~N524;
  assign T138 = ~N523;
  assign T140 = T142 & T141;
  assign T141 = ~sign_PA;
  assign T142 = T144 & T143;
  assign T143 = ~N519;
  assign T144 = ~N524;
  assign entering_PB = entering_PB_S | leaving_PA;
  assign entering_PB_S = T150 & T145;
  assign T145 = leaving_PB | T146;
  assign T146 = T148 & T147;
  assign T147 = ~ready_PC;
  assign T148 = ~valid_PB;
  assign leaving_PB = valid_PB & valid_leaving_PB;
  assign T150 = T152 & T151;
  assign T151 = ~valid_PA;
  assign T152 = cyc_S & T153;
  assign T153 = ~normalCase_S;
  assign T155 = entering_PB | leaving_PB;
  assign entering_PC = entering_PC_S | leaving_PB;
  assign entering_PC_S = T156 & ready_PC;
  assign T156 = T158 & T157;
  assign T157 = ~valid_PB;
  assign T158 = T160 & T159;
  assign T159 = ~valid_PA;
  assign T160 = cyc_S & T161;
  assign T161 = ~normalCase_S;
  assign N129 = ~T165;
  assign T163[53] = ~io_mulAddResult_3[104];
  assign T163[52] = ~io_mulAddResult_3[103];
  assign T163[51] = ~io_mulAddResult_3[102];
  assign T163[50] = ~io_mulAddResult_3[101];
  assign T163[49] = ~io_mulAddResult_3[100];
  assign T163[48] = ~io_mulAddResult_3[99];
  assign T163[47] = ~io_mulAddResult_3[98];
  assign T163[46] = ~io_mulAddResult_3[97];
  assign T163[45] = ~io_mulAddResult_3[96];
  assign T163[44] = ~io_mulAddResult_3[95];
  assign T163[43] = ~io_mulAddResult_3[94];
  assign T163[42] = ~io_mulAddResult_3[93];
  assign T163[41] = ~io_mulAddResult_3[92];
  assign T163[40] = ~io_mulAddResult_3[91];
  assign T163[39] = ~io_mulAddResult_3[90];
  assign T163[38] = ~io_mulAddResult_3[89];
  assign T163[37] = ~io_mulAddResult_3[88];
  assign T163[36] = ~io_mulAddResult_3[87];
  assign T163[35] = ~io_mulAddResult_3[86];
  assign T163[34] = ~io_mulAddResult_3[85];
  assign T163[33] = ~io_mulAddResult_3[84];
  assign T163[32] = ~io_mulAddResult_3[83];
  assign T163[31] = ~io_mulAddResult_3[82];
  assign T163[30] = ~io_mulAddResult_3[81];
  assign T163[29] = ~io_mulAddResult_3[80];
  assign T163[28] = ~io_mulAddResult_3[79];
  assign T163[27] = ~io_mulAddResult_3[78];
  assign T163[26] = ~io_mulAddResult_3[77];
  assign T163[25] = ~io_mulAddResult_3[76];
  assign T163[24] = ~io_mulAddResult_3[75];
  assign T163[23] = ~io_mulAddResult_3[74];
  assign T163[22] = ~io_mulAddResult_3[73];
  assign T163[21] = ~io_mulAddResult_3[72];
  assign T163[20] = ~io_mulAddResult_3[71];
  assign T163[19] = ~io_mulAddResult_3[70];
  assign T163[18] = ~io_mulAddResult_3[69];
  assign T163[17] = ~io_mulAddResult_3[68];
  assign T163[16] = ~io_mulAddResult_3[67];
  assign T163[15] = ~io_mulAddResult_3[66];
  assign T163[14] = ~io_mulAddResult_3[65];
  assign T163[13] = ~io_mulAddResult_3[64];
  assign T163[12] = ~io_mulAddResult_3[63];
  assign T163[11] = ~io_mulAddResult_3[62];
  assign T163[10] = ~io_mulAddResult_3[61];
  assign T163[9] = ~io_mulAddResult_3[60];
  assign T163[8] = ~io_mulAddResult_3[59];
  assign T163[7] = ~io_mulAddResult_3[58];
  assign T163[6] = ~io_mulAddResult_3[57];
  assign T163[5] = ~io_mulAddResult_3[56];
  assign T163[4] = ~io_mulAddResult_3[55];
  assign T163[3] = ~io_mulAddResult_3[54];
  assign T163[2] = ~io_mulAddResult_3[53];
  assign T163[1] = ~io_mulAddResult_3[52];
  assign T163[0] = ~io_mulAddResult_3[51];
  assign T165 = T166 | cyc_C1_sqrt;
  assign cyc_C1_sqrt = N312 & sqrtOp_PC;
  assign T166 = cyc_C1_div & T167;
  assign T167 = ~E_C1_div;
  assign N130 = ~exp_PC[0];
  assign entering_PB_normalCase = T177 & valid_normalCase_leaving_PA;
  assign T177 = valid_PA & normalCase_PA;
  assign entering_PC_normalCase = T178 & N509;
  assign T178 = valid_PB & normalCase_PB;
  assign T170[1] = sigB_PC[1] ^ T170[0];
  assign N131 = ~io_sqrtOp;
  assign T198[10] = ~io_b[62];
  assign T198[9] = ~io_b[61];
  assign T198[8] = ~io_b[60];
  assign T198[7] = ~io_b[59];
  assign T198[6] = ~io_b[58];
  assign T198[5] = ~io_b[57];
  assign T198[4] = ~io_b[56];
  assign T198[3] = ~io_b[55];
  assign T198[2] = ~io_b[54];
  assign T198[1] = ~io_b[53];
  assign T198[0] = ~io_b[52];
  assign cyc_E3_sqrt = N289 & sqrtOp_PC;
  assign T204[104] = T216[104] | 1'b0;
  assign T204[103] = T216[103] | 1'b0;
  assign T204[102] = T216[102] | 1'b0;
  assign T204[101] = T216[101] | 1'b0;
  assign T204[100] = T216[100] | 1'b0;
  assign T204[99] = T216[99] | 1'b0;
  assign T204[98] = T216[98] | 1'b0;
  assign T204[97] = T216[97] | 1'b0;
  assign T204[96] = T216[96] | 1'b0;
  assign T204[95] = T216[95] | 1'b0;
  assign T204[94] = T216[94] | 1'b0;
  assign T204[93] = T216[93] | 1'b0;
  assign T204[92] = T216[92] | 1'b0;
  assign T204[91] = T216[91] | 1'b0;
  assign T204[90] = T216[90] | 1'b0;
  assign T204[89] = T216[89] | 1'b0;
  assign T204[88] = T216[88] | 1'b0;
  assign T204[87] = T216[87] | 1'b0;
  assign T204[86] = T216[86] | 1'b0;
  assign T204[85] = T216[85] | 1'b0;
  assign T204[84] = T216[84] | 1'b0;
  assign T204[83] = T216[83] | 1'b0;
  assign T204[82] = T216[82] | 1'b0;
  assign T204[81] = T216[81] | 1'b0;
  assign T204[80] = T216[80] | 1'b0;
  assign T204[79] = T216[79] | 1'b0;
  assign T204[78] = T216[78] | 1'b0;
  assign T204[77] = T216[77] | 1'b0;
  assign T204[76] = T216[76] | 1'b0;
  assign T204[75] = T216[75] | 1'b0;
  assign T204[74] = T216[74] | 1'b0;
  assign T204[73] = T216[73] | 1'b0;
  assign T204[72] = T216[72] | 1'b0;
  assign T204[71] = T216[71] | 1'b0;
  assign T204[70] = T216[70] | 1'b0;
  assign T204[69] = T216[69] | 1'b0;
  assign T204[68] = T216[68] | 1'b0;
  assign T204[67] = T216[67] | 1'b0;
  assign T204[66] = T216[66] | 1'b0;
  assign T204[65] = T216[65] | 1'b0;
  assign T204[64] = T216[64] | 1'b0;
  assign T204[63] = T216[63] | 1'b0;
  assign T204[62] = T216[62] | 1'b0;
  assign T204[61] = T216[61] | 1'b0;
  assign T204[60] = T216[60] | 1'b0;
  assign T204[59] = T216[59] | 1'b0;
  assign T204[58] = T216[58] | 1'b0;
  assign T204[57] = T216[57] | 1'b0;
  assign T204[56] = T216[56] | 1'b0;
  assign T204[55] = T216[55] | 1'b0;
  assign T204[54] = T216[54] | 1'b0;
  assign T204[53] = T216[53] | T897[53];
  assign T204[52] = T216[52] | 1'b0;
  assign T204[51] = T216[51] | 1'b0;
  assign T204[50] = T216[50] | 1'b0;
  assign T204[49] = T216[49] | 1'b0;
  assign T204[48] = T216[48] | 1'b0;
  assign T204[47] = T216[47] | 1'b0;
  assign T204[46] = T216[46] | 1'b0;
  assign T204[45] = T216[45] | 1'b0;
  assign T204[44] = T216[44] | 1'b0;
  assign T204[43] = T216[43] | 1'b0;
  assign T204[42] = T216[42] | 1'b0;
  assign T204[41] = T216[41] | 1'b0;
  assign T204[40] = T216[40] | 1'b0;
  assign T204[39] = T216[39] | 1'b0;
  assign T204[38] = T216[38] | 1'b0;
  assign T204[37] = T216[37] | 1'b0;
  assign T204[36] = T216[36] | 1'b0;
  assign T204[35] = T216[35] | 1'b0;
  assign T204[34] = T216[34] | 1'b0;
  assign T204[33] = T216[33] | 1'b0;
  assign T204[32] = T216[32] | 1'b0;
  assign T204[31] = T216[31] | 1'b0;
  assign T204[30] = T216[30] | 1'b0;
  assign T204[29] = T216[29] | 1'b0;
  assign T204[28] = T216[28] | 1'b0;
  assign T204[27] = T216[27] | 1'b0;
  assign T204[26] = T216[26] | 1'b0;
  assign T204[25] = T216[25] | 1'b0;
  assign T204[24] = T216[24] | 1'b0;
  assign T204[23] = T216[23] | 1'b0;
  assign T204[22] = T216[22] | 1'b0;
  assign T204[21] = T216[21] | 1'b0;
  assign T204[20] = T216[20] | 1'b0;
  assign T204[19] = T216[19] | 1'b0;
  assign T204[18] = T216[18] | 1'b0;
  assign T204[17] = T216[17] | 1'b0;
  assign T204[16] = T216[16] | 1'b0;
  assign T204[15] = T216[15] | 1'b0;
  assign T204[14] = T216[14] | 1'b0;
  assign T204[13] = T216[13] | 1'b0;
  assign T204[12] = T216[12] | 1'b0;
  assign T204[11] = T216[11] | 1'b0;
  assign T204[10] = T216[10] | 1'b0;
  assign T204[9] = T216[9] | 1'b0;
  assign T204[8] = T216[8] | 1'b0;
  assign T204[7] = T216[7] | 1'b0;
  assign T204[6] = T216[6] | 1'b0;
  assign T204[5] = T216[5] | 1'b0;
  assign T204[4] = T216[4] | 1'b0;
  assign T204[3] = T216[3] | 1'b0;
  assign T204[2] = T216[2] | 1'b0;
  assign T204[1] = T216[1] | 1'b0;
  assign T204[0] = T216[0] | 1'b0;
  assign N132 = ~T212;
  assign T212 = cyc_E3_div & T213;
  assign T213 = ~E_E_div;
  assign cyc_E3_div = N289 & T215;
  assign T215 = ~sqrtOp_PC;
  assign T216[104] = T228[104] | T217[104];
  assign T216[103] = T228[103] | T217[103];
  assign T216[102] = T228[102] | T217[102];
  assign T216[101] = T228[101] | T217[101];
  assign T216[100] = T228[100] | T217[100];
  assign T216[99] = T228[99] | T217[99];
  assign T216[98] = T228[98] | T217[98];
  assign T216[97] = T228[97] | T217[97];
  assign T216[96] = T228[96] | T217[96];
  assign T216[95] = T228[95] | T217[95];
  assign T216[94] = T228[94] | T217[94];
  assign T216[93] = T228[93] | T217[93];
  assign T216[92] = T228[92] | T217[92];
  assign T216[91] = T228[91] | T217[91];
  assign T216[90] = T228[90] | T217[90];
  assign T216[89] = T228[89] | T217[89];
  assign T216[88] = T228[88] | T217[88];
  assign T216[87] = T228[87] | T217[87];
  assign T216[86] = T228[86] | T217[86];
  assign T216[85] = T228[85] | T217[85];
  assign T216[84] = T228[84] | T217[84];
  assign T216[83] = T228[83] | T217[83];
  assign T216[82] = T228[82] | T217[82];
  assign T216[81] = T228[81] | T217[81];
  assign T216[80] = T228[80] | T217[80];
  assign T216[79] = T228[79] | T217[79];
  assign T216[78] = T228[78] | T217[78];
  assign T216[77] = T228[77] | T217[77];
  assign T216[76] = T228[76] | T217[76];
  assign T216[75] = T228[75] | T217[75];
  assign T216[74] = T228[74] | T217[74];
  assign T216[73] = T228[73] | T217[73];
  assign T216[72] = T228[72] | T217[72];
  assign T216[71] = T228[71] | T217[71];
  assign T216[70] = T228[70] | T217[70];
  assign T216[69] = T228[69] | T217[69];
  assign T216[68] = T228[68] | T217[68];
  assign T216[67] = T228[67] | T217[67];
  assign T216[66] = T228[66] | T217[66];
  assign T216[65] = T228[65] | T217[65];
  assign T216[64] = T228[64] | T217[64];
  assign T216[63] = T228[63] | T217[63];
  assign T216[62] = T228[62] | T217[62];
  assign T216[61] = T228[61] | T217[61];
  assign T216[60] = T228[60] | T217[60];
  assign T216[59] = T228[59] | T217[59];
  assign T216[58] = T228[58] | T217[58];
  assign T216[57] = T228[57] | T217[57];
  assign T216[56] = T228[56] | T217[56];
  assign T216[55] = T228[55] | T217[55];
  assign T216[54] = T228[54] | T217[54];
  assign T216[53] = T228[53] | T217[53];
  assign T216[52] = T228[52] | T217[52];
  assign T216[51] = T228[51] | T217[51];
  assign T216[50] = T228[50] | T217[50];
  assign T216[49] = T228[49] | T217[49];
  assign T216[48] = T228[48] | T217[48];
  assign T216[47] = T228[47] | T217[47];
  assign T216[46] = T228[46] | 1'b0;
  assign T216[45] = T228[45] | 1'b0;
  assign T216[44] = T228[44] | 1'b0;
  assign T216[43] = T228[43] | 1'b0;
  assign T216[42] = T228[42] | 1'b0;
  assign T216[41] = T228[41] | 1'b0;
  assign T216[40] = T228[40] | 1'b0;
  assign T216[39] = T228[39] | 1'b0;
  assign T216[38] = T228[38] | 1'b0;
  assign T216[37] = T228[37] | 1'b0;
  assign T216[36] = T228[36] | 1'b0;
  assign T216[35] = T228[35] | 1'b0;
  assign T216[34] = T228[34] | 1'b0;
  assign T216[33] = T228[33] | 1'b0;
  assign T216[32] = T228[32] | 1'b0;
  assign T216[31] = T228[31] | 1'b0;
  assign T216[30] = T228[30] | 1'b0;
  assign T216[29] = T228[29] | 1'b0;
  assign T216[28] = T228[28] | 1'b0;
  assign T216[27] = T228[27] | 1'b0;
  assign T216[26] = T228[26] | 1'b0;
  assign T216[25] = T228[25] | 1'b0;
  assign T216[24] = T228[24] | 1'b0;
  assign T216[23] = T228[23] | 1'b0;
  assign T216[22] = T228[22] | 1'b0;
  assign T216[21] = T228[21] | 1'b0;
  assign T216[20] = T228[20] | 1'b0;
  assign T216[19] = T228[19] | 1'b0;
  assign T216[18] = T228[18] | 1'b0;
  assign T216[17] = T228[17] | 1'b0;
  assign T216[16] = T228[16] | 1'b0;
  assign T216[15] = T228[15] | 1'b0;
  assign T216[14] = T228[14] | 1'b0;
  assign T216[13] = T228[13] | 1'b0;
  assign T216[12] = T228[12] | 1'b0;
  assign T216[11] = T228[11] | 1'b0;
  assign T216[10] = T228[10] | 1'b0;
  assign T216[9] = T228[9] | 1'b0;
  assign T216[8] = T228[8] | 1'b0;
  assign T216[7] = T228[7] | 1'b0;
  assign T216[6] = T228[6] | 1'b0;
  assign T216[5] = T228[5] | 1'b0;
  assign T216[4] = T228[4] | 1'b0;
  assign T216[3] = T228[3] | 1'b0;
  assign T216[2] = T228[2] | 1'b0;
  assign T216[1] = T228[1] | 1'b0;
  assign T216[0] = T228[0] | 1'b0;
  assign N133 = ~T225;
  assign T221 = T222 | cyc_C3_sqrt;
  assign cyc_C3_sqrt = N509 & sqrtOp_PB;
  assign T222 = N308 | cyc_C5_div;
  assign cyc_C5_div = N481 & T223;
  assign T223 = ~sqrtOp_PB;
  assign T225 = cyc_C4_sqrt | N285;
  assign cyc_C4_sqrt = N476 & sqrtOp_PB;
  assign T228[104] = T233[104] | 1'b0;
  assign T228[103] = T233[103] | T898[103];
  assign T228[102] = T233[102] | T898[102];
  assign T228[101] = T233[101] | T898[101];
  assign T228[100] = T233[100] | T898[100];
  assign T228[99] = T233[99] | T898[99];
  assign T228[98] = T233[98] | T898[98];
  assign T228[97] = T233[97] | T898[97];
  assign T228[96] = T233[96] | T898[96];
  assign T228[95] = T233[95] | T898[95];
  assign T228[94] = T233[94] | T898[94];
  assign T228[93] = T233[93] | T898[93];
  assign T228[92] = T233[92] | T898[92];
  assign T228[91] = T233[91] | T898[91];
  assign T228[90] = T233[90] | T898[90];
  assign T228[89] = T233[89] | T898[89];
  assign T228[88] = T233[88] | T898[88];
  assign T228[87] = T233[87] | T898[87];
  assign T228[86] = T233[86] | T898[86];
  assign T228[85] = T233[85] | T898[85];
  assign T228[84] = T233[84] | T898[84];
  assign T228[83] = T233[83] | T898[83];
  assign T228[82] = T233[82] | T898[82];
  assign T228[81] = T233[81] | T898[81];
  assign T228[80] = T233[80] | T898[80];
  assign T228[79] = T233[79] | T898[79];
  assign T228[78] = T233[78] | T898[78];
  assign T228[77] = T233[77] | T898[77];
  assign T228[76] = T233[76] | T898[76];
  assign T228[75] = T233[75] | T898[75];
  assign T228[74] = T233[74] | T898[74];
  assign T228[73] = T233[73] | T898[73];
  assign T228[72] = T233[72] | T898[72];
  assign T228[71] = T233[71] | T898[71];
  assign T228[70] = T233[70] | T898[70];
  assign T228[69] = T233[69] | T898[69];
  assign T228[68] = T233[68] | T898[68];
  assign T228[67] = T233[67] | T898[67];
  assign T228[66] = T233[66] | T898[66];
  assign T228[65] = T233[65] | T898[65];
  assign T228[64] = T233[64] | T898[64];
  assign T228[63] = T233[63] | T898[63];
  assign T228[62] = T233[62] | T898[62];
  assign T228[61] = T233[61] | T898[61];
  assign T228[60] = T233[60] | T898[60];
  assign T228[59] = T233[59] | T898[59];
  assign T228[58] = T233[58] | T898[58];
  assign T228[57] = T233[57] | T898[57];
  assign T228[56] = T233[56] | T898[56];
  assign T228[55] = T233[55] | T898[55];
  assign T228[54] = T233[54] | T898[54];
  assign T228[53] = T233[53] | T898[53];
  assign T228[52] = T233[52] | T898[52];
  assign T228[51] = T233[51] | T898[51];
  assign T228[50] = T233[50] | T898[50];
  assign T228[49] = T233[49] | T898[49];
  assign T228[48] = T233[48] | T898[48];
  assign T228[47] = T233[47] | T898[47];
  assign T228[46] = 1'b0 | T898[46];
  assign T228[45] = 1'b0 | 1'b0;
  assign T228[44] = 1'b0 | 1'b0;
  assign T228[43] = 1'b0 | 1'b0;
  assign T228[42] = 1'b0 | 1'b0;
  assign T228[41] = 1'b0 | 1'b0;
  assign T228[40] = 1'b0 | 1'b0;
  assign T228[39] = 1'b0 | 1'b0;
  assign T228[38] = 1'b0 | 1'b0;
  assign T228[37] = 1'b0 | 1'b0;
  assign T228[36] = 1'b0 | 1'b0;
  assign T228[35] = 1'b0 | 1'b0;
  assign T228[34] = 1'b0 | 1'b0;
  assign T228[33] = 1'b0 | 1'b0;
  assign T228[32] = 1'b0 | 1'b0;
  assign T228[31] = 1'b0 | 1'b0;
  assign T228[30] = 1'b0 | 1'b0;
  assign T228[29] = 1'b0 | 1'b0;
  assign T228[28] = 1'b0 | 1'b0;
  assign T228[27] = 1'b0 | 1'b0;
  assign T228[26] = 1'b0 | 1'b0;
  assign T228[25] = 1'b0 | 1'b0;
  assign T228[24] = 1'b0 | 1'b0;
  assign T228[23] = 1'b0 | 1'b0;
  assign T228[22] = 1'b0 | 1'b0;
  assign T228[21] = 1'b0 | 1'b0;
  assign T228[20] = 1'b0 | 1'b0;
  assign T228[19] = 1'b0 | 1'b0;
  assign T228[18] = 1'b0 | 1'b0;
  assign T228[17] = 1'b0 | 1'b0;
  assign T228[16] = 1'b0 | 1'b0;
  assign T228[15] = 1'b0 | 1'b0;
  assign T228[14] = 1'b0 | 1'b0;
  assign T228[13] = 1'b0 | 1'b0;
  assign T228[12] = 1'b0 | 1'b0;
  assign T228[11] = 1'b0 | 1'b0;
  assign T228[10] = 1'b0 | 1'b0;
  assign T228[9] = 1'b0 | 1'b0;
  assign T228[8] = 1'b0 | 1'b0;
  assign T228[7] = 1'b0 | 1'b0;
  assign T228[6] = 1'b0 | 1'b0;
  assign T228[5] = 1'b0 | 1'b0;
  assign T228[4] = 1'b0 | 1'b0;
  assign T228[3] = 1'b0 | 1'b0;
  assign T228[2] = 1'b0 | 1'b0;
  assign T228[1] = 1'b0 | 1'b0;
  assign T228[0] = 1'b0 | 1'b0;
  assign io_mulAddB_0[53] = 1'b0 | zComplSigT_C1[53];
  assign io_mulAddB_0[52] = T899[52] | zComplSigT_C1[52];
  assign io_mulAddB_0[51] = T899[51] | zComplSigT_C1[51];
  assign io_mulAddB_0[50] = T899[50] | zComplSigT_C1[50];
  assign io_mulAddB_0[49] = T899[49] | zComplSigT_C1[49];
  assign io_mulAddB_0[48] = T899[48] | zComplSigT_C1[48];
  assign io_mulAddB_0[47] = T899[47] | zComplSigT_C1[47];
  assign io_mulAddB_0[46] = T899[46] | zComplSigT_C1[46];
  assign io_mulAddB_0[45] = T899[45] | zComplSigT_C1[45];
  assign io_mulAddB_0[44] = T899[44] | zComplSigT_C1[44];
  assign io_mulAddB_0[43] = T899[43] | zComplSigT_C1[43];
  assign io_mulAddB_0[42] = T899[42] | zComplSigT_C1[42];
  assign io_mulAddB_0[41] = T899[41] | zComplSigT_C1[41];
  assign io_mulAddB_0[40] = T899[40] | zComplSigT_C1[40];
  assign io_mulAddB_0[39] = T899[39] | zComplSigT_C1[39];
  assign io_mulAddB_0[38] = T899[38] | zComplSigT_C1[38];
  assign io_mulAddB_0[37] = T899[37] | zComplSigT_C1[37];
  assign io_mulAddB_0[36] = T899[36] | zComplSigT_C1[36];
  assign io_mulAddB_0[35] = T899[35] | zComplSigT_C1[35];
  assign io_mulAddB_0[34] = T899[34] | zComplSigT_C1[34];
  assign io_mulAddB_0[33] = T899[33] | zComplSigT_C1[33];
  assign io_mulAddB_0[32] = T899[32] | zComplSigT_C1[32];
  assign io_mulAddB_0[31] = T899[31] | zComplSigT_C1[31];
  assign io_mulAddB_0[30] = T899[30] | zComplSigT_C1[30];
  assign io_mulAddB_0[29] = T899[29] | zComplSigT_C1[29];
  assign io_mulAddB_0[28] = T899[28] | zComplSigT_C1[28];
  assign io_mulAddB_0[27] = T899[27] | zComplSigT_C1[27];
  assign io_mulAddB_0[26] = T899[26] | zComplSigT_C1[26];
  assign io_mulAddB_0[25] = T899[25] | zComplSigT_C1[25];
  assign io_mulAddB_0[24] = T899[24] | zComplSigT_C1[24];
  assign io_mulAddB_0[23] = T899[23] | zComplSigT_C1[23];
  assign io_mulAddB_0[22] = T899[22] | zComplSigT_C1[22];
  assign io_mulAddB_0[21] = T899[21] | zComplSigT_C1[21];
  assign io_mulAddB_0[20] = T899[20] | zComplSigT_C1[20];
  assign io_mulAddB_0[19] = T899[19] | zComplSigT_C1[19];
  assign io_mulAddB_0[18] = T899[18] | zComplSigT_C1[18];
  assign io_mulAddB_0[17] = T899[17] | zComplSigT_C1[17];
  assign io_mulAddB_0[16] = T899[16] | zComplSigT_C1[16];
  assign io_mulAddB_0[15] = T899[15] | zComplSigT_C1[15];
  assign io_mulAddB_0[14] = T899[14] | zComplSigT_C1[14];
  assign io_mulAddB_0[13] = T899[13] | zComplSigT_C1[13];
  assign io_mulAddB_0[12] = T899[12] | zComplSigT_C1[12];
  assign io_mulAddB_0[11] = T899[11] | zComplSigT_C1[11];
  assign io_mulAddB_0[10] = T899[10] | zComplSigT_C1[10];
  assign io_mulAddB_0[9] = T899[9] | zComplSigT_C1[9];
  assign io_mulAddB_0[8] = T899[8] | zComplSigT_C1[8];
  assign io_mulAddB_0[7] = T899[7] | zComplSigT_C1[7];
  assign io_mulAddB_0[6] = T899[6] | zComplSigT_C1[6];
  assign io_mulAddB_0[5] = T899[5] | zComplSigT_C1[5];
  assign io_mulAddB_0[4] = T899[4] | zComplSigT_C1[4];
  assign io_mulAddB_0[3] = T899[3] | zComplSigT_C1[3];
  assign io_mulAddB_0[2] = T899[2] | zComplSigT_C1[2];
  assign io_mulAddB_0[1] = T899[1] | zComplSigT_C1[1];
  assign io_mulAddB_0[0] = T899[0] | zComplSigT_C1[0];
  assign T899[52] = T239[52] | 1'b0;
  assign T899[51] = T239[51] | 1'b0;
  assign T899[50] = T239[50] | 1'b0;
  assign T899[49] = T239[49] | 1'b0;
  assign T899[48] = T239[48] | 1'b0;
  assign T899[47] = T239[47] | 1'b0;
  assign T899[46] = T239[46] | 1'b0;
  assign T899[45] = T239[45] | 1'b0;
  assign T899[44] = T239[44] | 1'b0;
  assign T899[43] = T239[43] | 1'b0;
  assign T899[42] = T239[42] | 1'b0;
  assign T899[41] = T239[41] | 1'b0;
  assign T899[40] = T239[40] | 1'b0;
  assign T899[39] = T239[39] | 1'b0;
  assign T899[38] = T239[38] | 1'b0;
  assign T899[37] = T239[37] | 1'b0;
  assign T899[36] = T239[36] | 1'b0;
  assign T899[35] = T239[35] | 1'b0;
  assign T899[34] = T239[34] | 1'b0;
  assign T899[33] = T239[33] | 1'b0;
  assign T899[32] = T239[32] | T900[32];
  assign T899[31] = T239[31] | T900[31];
  assign T899[30] = T239[30] | T900[30];
  assign T899[29] = T239[29] | T900[29];
  assign T899[28] = T239[28] | T900[28];
  assign T899[27] = T239[27] | T900[27];
  assign T899[26] = T239[26] | T900[26];
  assign T899[25] = T239[25] | T900[25];
  assign T899[24] = T239[24] | T900[24];
  assign T899[23] = T239[23] | T900[23];
  assign T899[22] = T239[22] | T900[22];
  assign T899[21] = T239[21] | T900[21];
  assign T899[20] = T239[20] | T900[20];
  assign T899[19] = T239[19] | T900[19];
  assign T899[18] = T239[18] | T900[18];
  assign T899[17] = T239[17] | T900[17];
  assign T899[16] = T239[16] | T900[16];
  assign T899[15] = T239[15] | T900[15];
  assign T899[14] = T239[14] | T900[14];
  assign T899[13] = T239[13] | T900[13];
  assign T899[12] = T239[12] | T900[12];
  assign T899[11] = T239[11] | T900[11];
  assign T899[10] = T239[10] | T900[10];
  assign T899[9] = T239[9] | T900[9];
  assign T899[8] = T239[8] | T900[8];
  assign T899[7] = T239[7] | T900[7];
  assign T899[6] = T239[6] | T900[6];
  assign T899[5] = T239[5] | T900[5];
  assign T899[4] = T239[4] | T900[4];
  assign T899[3] = T239[3] | T900[3];
  assign T899[2] = T239[2] | T900[2];
  assign T899[1] = T239[1] | T900[1];
  assign T899[0] = T239[0] | T900[0];
  assign T239[52] = T242[52] | 1'b0;
  assign T239[51] = T242[51] | 1'b0;
  assign T239[50] = T242[50] | 1'b0;
  assign T239[49] = T242[49] | 1'b0;
  assign T239[48] = T242[48] | 1'b0;
  assign T239[47] = T242[47] | 1'b0;
  assign T239[46] = T242[46] | 1'b0;
  assign T239[45] = T242[45] | 1'b0;
  assign T239[44] = T242[44] | 1'b0;
  assign T239[43] = T242[43] | 1'b0;
  assign T239[42] = T242[42] | 1'b0;
  assign T239[41] = T242[41] | 1'b0;
  assign T239[40] = T242[40] | 1'b0;
  assign T239[39] = T242[39] | 1'b0;
  assign T239[38] = T242[38] | 1'b0;
  assign T239[37] = T242[37] | 1'b0;
  assign T239[36] = T242[36] | 1'b0;
  assign T239[35] = T242[35] | 1'b0;
  assign T239[34] = T242[34] | 1'b0;
  assign T239[33] = T242[33] | 1'b0;
  assign T239[32] = T242[32] | 1'b0;
  assign T239[31] = T242[31] | 1'b0;
  assign T239[30] = T242[30] | 1'b0;
  assign T239[29] = T242[29] | T901[29];
  assign T239[28] = T242[28] | T901[28];
  assign T239[27] = T242[27] | T901[27];
  assign T239[26] = T242[26] | T901[26];
  assign T239[25] = T242[25] | T901[25];
  assign T239[24] = T242[24] | T901[24];
  assign T239[23] = T242[23] | T901[23];
  assign T239[22] = T242[22] | T901[22];
  assign T239[21] = T242[21] | T901[21];
  assign T239[20] = T242[20] | T901[20];
  assign T239[19] = T242[19] | T901[19];
  assign T239[18] = T242[18] | T901[18];
  assign T239[17] = T242[17] | T901[17];
  assign T239[16] = T242[16] | T901[16];
  assign T239[15] = T242[15] | T901[15];
  assign T239[14] = T242[14] | T901[14];
  assign T239[13] = T242[13] | T901[13];
  assign T239[12] = T242[12] | T901[12];
  assign T239[11] = T242[11] | T901[11];
  assign T239[10] = T242[10] | T901[10];
  assign T239[9] = T242[9] | T901[9];
  assign T239[8] = T242[8] | T901[8];
  assign T239[7] = T242[7] | T901[7];
  assign T239[6] = T242[6] | T901[6];
  assign T239[5] = T242[5] | T901[5];
  assign T239[4] = T242[4] | T901[4];
  assign T239[3] = T242[3] | T901[3];
  assign T239[2] = T242[2] | T901[2];
  assign T239[1] = T242[1] | T901[1];
  assign T239[0] = T242[0] | T901[0];
  assign T242[52] = T246[52] | 1'b0;
  assign T242[51] = T246[51] | 1'b0;
  assign T242[50] = T246[50] | 1'b0;
  assign T242[49] = T246[49] | 1'b0;
  assign T242[48] = T246[48] | 1'b0;
  assign T242[47] = T246[47] | 1'b0;
  assign T242[46] = T246[46] | 1'b0;
  assign T242[45] = T246[45] | T902[45];
  assign T242[44] = T246[44] | T902[44];
  assign T242[43] = T246[43] | T902[43];
  assign T242[42] = T246[42] | T902[42];
  assign T242[41] = T246[41] | T902[41];
  assign T242[40] = T246[40] | T902[40];
  assign T242[39] = T246[39] | T902[39];
  assign T242[38] = T246[38] | T902[38];
  assign T242[37] = T246[37] | T902[37];
  assign T242[36] = T246[36] | T902[36];
  assign T242[35] = T246[35] | T902[35];
  assign T242[34] = T246[34] | T902[34];
  assign T242[33] = T246[33] | T902[33];
  assign T242[32] = T246[32] | T902[32];
  assign T242[31] = T246[31] | T902[31];
  assign T242[30] = T246[30] | T902[30];
  assign T242[29] = T246[29] | T902[29];
  assign T242[28] = T246[28] | T902[28];
  assign T242[27] = T246[27] | T902[27];
  assign T242[26] = T246[26] | T902[26];
  assign T242[25] = T246[25] | T902[25];
  assign T242[24] = T246[24] | T902[24];
  assign T242[23] = T246[23] | T902[23];
  assign T242[22] = T246[22] | T902[22];
  assign T242[21] = T246[21] | T902[21];
  assign T242[20] = T246[20] | T902[20];
  assign T242[19] = T246[19] | T902[19];
  assign T242[18] = T246[18] | T902[18];
  assign T242[17] = T246[17] | T902[17];
  assign T242[16] = T246[16] | T902[16];
  assign T242[15] = T246[15] | T902[15];
  assign T242[14] = T246[14] | T902[14];
  assign T242[13] = T246[13] | T902[13];
  assign T242[12] = T246[12] | T902[12];
  assign T242[11] = T246[11] | T902[11];
  assign T242[10] = T246[10] | T902[10];
  assign T242[9] = T246[9] | T902[9];
  assign T242[8] = T246[8] | T902[8];
  assign T242[7] = T246[7] | T902[7];
  assign T242[6] = T246[6] | T902[6];
  assign T242[5] = T246[5] | T902[5];
  assign T242[4] = T246[4] | T902[4];
  assign T242[3] = T246[3] | T902[3];
  assign T242[2] = T246[2] | T902[2];
  assign T242[1] = T246[1] | T902[1];
  assign T242[0] = T246[0] | T902[0];
  assign T244[45] = ~io_mulAddResult_3[90];
  assign T244[44] = ~io_mulAddResult_3[89];
  assign T244[43] = ~io_mulAddResult_3[88];
  assign T244[42] = ~io_mulAddResult_3[87];
  assign T244[41] = ~io_mulAddResult_3[86];
  assign T244[40] = ~io_mulAddResult_3[85];
  assign T244[39] = ~io_mulAddResult_3[84];
  assign T244[38] = ~io_mulAddResult_3[83];
  assign T244[37] = ~io_mulAddResult_3[82];
  assign T244[36] = ~io_mulAddResult_3[81];
  assign T244[35] = ~io_mulAddResult_3[80];
  assign T244[34] = ~io_mulAddResult_3[79];
  assign T244[33] = ~io_mulAddResult_3[78];
  assign T244[32] = ~io_mulAddResult_3[77];
  assign T244[31] = ~io_mulAddResult_3[76];
  assign T244[30] = ~io_mulAddResult_3[75];
  assign T244[29] = ~io_mulAddResult_3[74];
  assign T244[28] = ~io_mulAddResult_3[73];
  assign T244[27] = ~io_mulAddResult_3[72];
  assign T244[26] = ~io_mulAddResult_3[71];
  assign T244[25] = ~io_mulAddResult_3[70];
  assign T244[24] = ~io_mulAddResult_3[69];
  assign T244[23] = ~io_mulAddResult_3[68];
  assign T244[22] = ~io_mulAddResult_3[67];
  assign T244[21] = ~io_mulAddResult_3[66];
  assign T244[20] = ~io_mulAddResult_3[65];
  assign T244[19] = ~io_mulAddResult_3[64];
  assign T244[18] = ~io_mulAddResult_3[63];
  assign T244[17] = ~io_mulAddResult_3[62];
  assign T244[16] = ~io_mulAddResult_3[61];
  assign T244[15] = ~io_mulAddResult_3[60];
  assign T244[14] = ~io_mulAddResult_3[59];
  assign T244[13] = ~io_mulAddResult_3[58];
  assign T244[12] = ~io_mulAddResult_3[57];
  assign T244[11] = ~io_mulAddResult_3[56];
  assign T244[10] = ~io_mulAddResult_3[55];
  assign T244[9] = ~io_mulAddResult_3[54];
  assign T244[8] = ~io_mulAddResult_3[53];
  assign T244[7] = ~io_mulAddResult_3[52];
  assign T244[6] = ~io_mulAddResult_3[51];
  assign T244[5] = ~io_mulAddResult_3[50];
  assign T244[4] = ~io_mulAddResult_3[49];
  assign T244[3] = ~io_mulAddResult_3[48];
  assign T244[2] = ~io_mulAddResult_3[47];
  assign T244[1] = ~io_mulAddResult_3[46];
  assign T244[0] = ~io_mulAddResult_3[45];
  assign T246[52] = 1'b0 | T247[52];
  assign T246[51] = T925[51] | T247[51];
  assign T246[50] = T925[50] | T247[50];
  assign T246[49] = T925[49] | T247[49];
  assign T246[48] = T925[48] | T247[48];
  assign T246[47] = T925[47] | T247[47];
  assign T246[46] = T925[46] | T247[46];
  assign T246[45] = T925[45] | T247[45];
  assign T246[44] = T925[44] | T247[44];
  assign T246[43] = T925[43] | T247[43];
  assign T246[42] = T925[42] | T247[42];
  assign T246[41] = T925[41] | T247[41];
  assign T246[40] = T925[40] | T247[40];
  assign T246[39] = T925[39] | T247[39];
  assign T246[38] = T925[38] | T247[38];
  assign T246[37] = T925[37] | T247[37];
  assign T246[36] = T925[36] | T247[36];
  assign T246[35] = T925[35] | 1'b0;
  assign T246[34] = T925[34] | 1'b0;
  assign T246[33] = T925[33] | 1'b0;
  assign T246[32] = T925[32] | 1'b0;
  assign T246[31] = T925[31] | 1'b0;
  assign T246[30] = T925[30] | 1'b0;
  assign T246[29] = T925[29] | 1'b0;
  assign T246[28] = T925[28] | 1'b0;
  assign T246[27] = T925[27] | 1'b0;
  assign T246[26] = T925[26] | 1'b0;
  assign T246[25] = T925[25] | 1'b0;
  assign T246[24] = T925[24] | 1'b0;
  assign T246[23] = T925[23] | 1'b0;
  assign T246[22] = T925[22] | 1'b0;
  assign T246[21] = T925[21] | 1'b0;
  assign T246[20] = T925[20] | 1'b0;
  assign T246[19] = T925[19] | 1'b0;
  assign T246[18] = T925[18] | 1'b0;
  assign T246[17] = T925[17] | 1'b0;
  assign T246[16] = T925[16] | 1'b0;
  assign T246[15] = T925[15] | 1'b0;
  assign T246[14] = T925[14] | 1'b0;
  assign T246[13] = T925[13] | 1'b0;
  assign T246[12] = T925[12] | 1'b0;
  assign T246[11] = T925[11] | 1'b0;
  assign T246[10] = T925[10] | 1'b0;
  assign T246[9] = T925[9] | 1'b0;
  assign T246[8] = T925[8] | 1'b0;
  assign T246[7] = T925[7] | 1'b0;
  assign T246[6] = T925[6] | 1'b0;
  assign T246[5] = T925[5] | 1'b0;
  assign T246[4] = T925[4] | 1'b0;
  assign T246[3] = T925[3] | 1'b0;
  assign T246[2] = T925[2] | 1'b0;
  assign T246[1] = T925[1] | 1'b0;
  assign T246[0] = T925[0] | 1'b0;
  assign N134 = ~cyc_B6_sqrt;
  assign N135 = ~exp_PA[0];
  assign ER1_A1_sqrt[16] = exp_PA[0];
  assign mulAdd9C_A[24] = T271[24] | 1'b0;
  assign mulAdd9C_A[23] = T271[23] | T904[23];
  assign mulAdd9C_A[22] = T271[22] | T904[22];
  assign mulAdd9C_A[21] = T271[21] | T904[21];
  assign mulAdd9C_A[20] = T271[20] | T904[20];
  assign mulAdd9C_A[19] = T271[19] | T904[19];
  assign mulAdd9C_A[18] = T271[18] | T904[18];
  assign T253[17] = T271[17] | T904[17];
  assign T253[16] = T271[16] | T904[16];
  assign T253[15] = T271[15] | T904[15];
  assign T253[14] = T271[14] | 1'b0;
  assign T253[13] = T271[13] | 1'b0;
  assign T253[12] = T271[12] | 1'b0;
  assign T253[11] = T271[11] | 1'b0;
  assign T253[10] = T271[10] | 1'b0;
  assign T253[9] = T271[9] | 1'b0;
  assign T253[8] = T271[8] | 1'b0;
  assign T253[7] = T271[7] | 1'b0;
  assign T253[6] = T271[6] | 1'b0;
  assign T253[5] = T271[5] | 1'b0;
  assign T253[4] = T271[4] | 1'b0;
  assign T253[3] = T271[3] | 1'b0;
  assign T253[2] = T271[2] | 1'b0;
  assign T253[1] = T271[1] | 1'b0;
  assign T253[0] = T271[0] | 1'b0;
  assign N136 = ~cyc_A1_div;
  assign T258[8] = zFractR0_A6_sqrt[8] | zFractR0_A4_div[8];
  assign T258[7] = zFractR0_A6_sqrt[7] | zFractR0_A4_div[7];
  assign T258[6] = zFractR0_A6_sqrt[6] | zFractR0_A4_div[6];
  assign T258[5] = zFractR0_A6_sqrt[5] | zFractR0_A4_div[5];
  assign T258[4] = zFractR0_A6_sqrt[4] | zFractR0_A4_div[4];
  assign T258[3] = zFractR0_A6_sqrt[3] | zFractR0_A4_div[3];
  assign T258[2] = zFractR0_A6_sqrt[2] | zFractR0_A4_div[2];
  assign T258[1] = zFractR0_A6_sqrt[1] | zFractR0_A4_div[1];
  assign T258[0] = zFractR0_A6_sqrt[0] | zFractR0_A4_div[0];
  assign N137 = ~T262;
  assign T260[8] = ~T251[10];
  assign T260[7] = ~T251[9];
  assign T260[6] = ~T251[8];
  assign T260[5] = ~T251[7];
  assign T260[4] = ~T251[6];
  assign T260[3] = ~T251[5];
  assign T260[2] = ~T251[4];
  assign T260[1] = ~T251[3];
  assign T260[0] = ~T251[2];
  assign T262 = T305[20] & T251[11];
  assign N138 = ~T267;
  assign T265[8] = ~T251[9];
  assign T265[7] = ~T251[8];
  assign T265[6] = ~T251[7];
  assign T265[5] = ~T251[6];
  assign T265[4] = ~T251[5];
  assign T265[3] = ~T251[4];
  assign T265[2] = ~T251[3];
  assign T265[1] = ~T251[2];
  assign T265[0] = ~T251[1];
  assign T267 = N349 & T251[10];
  assign T269 = N349 | T305[20];
  assign cyc_A1_div = N316 & T270;
  assign T270 = ~sqrtOp_PA;
  assign T271[24] = 1'b0 | T272[24];
  assign T271[23] = 1'b0 | T272[23];
  assign T271[22] = 1'b0 | T272[22];
  assign T271[21] = 1'b0 | T272[21];
  assign T271[20] = T905[20] | T272[20];
  assign T271[19] = T905[19] | T272[19];
  assign T271[18] = T905[18] | T272[18];
  assign T271[17] = T905[17] | T272[17];
  assign T271[16] = T905[16] | T272[16];
  assign T271[15] = T905[15] | 1'b0;
  assign T271[14] = T905[14] | 1'b0;
  assign T271[13] = T905[13] | 1'b0;
  assign T271[12] = T905[12] | 1'b0;
  assign T271[11] = T905[11] | 1'b0;
  assign T271[10] = T905[10] | 1'b0;
  assign T271[9] = T905[9] | 1'b0;
  assign T271[8] = T905[8] | 1'b0;
  assign T271[7] = T905[7] | 1'b0;
  assign T271[6] = T905[6] | 1'b0;
  assign T271[5] = T905[5] | 1'b0;
  assign T271[4] = T905[4] | 1'b0;
  assign T271[3] = T905[3] | 1'b0;
  assign T271[2] = T905[2] | 1'b0;
  assign T271[1] = T905[1] | 1'b0;
  assign T271[0] = T905[0] | 1'b0;
  assign N139 = ~cyc_A1_sqrt;
  assign T905[20] = T282[20] | T275[20];
  assign T905[19] = T282[19] | T275[19];
  assign T905[18] = T282[18] | T275[18];
  assign T905[17] = T282[17] | T275[17];
  assign T905[16] = T282[16] | T275[16];
  assign T905[15] = T282[15] | T275[15];
  assign T905[14] = T282[14] | T275[14];
  assign T905[13] = T282[13] | T275[13];
  assign T905[12] = T282[12] | T275[12];
  assign T905[11] = T282[11] | T275[11];
  assign T905[10] = T282[10] | T275[10];
  assign T905[9] = T282[9] | T275[9];
  assign T905[8] = T282[8] | T275[8];
  assign T905[7] = T282[7] | T275[7];
  assign T905[6] = T282[6] | T275[6];
  assign T905[5] = T282[5] | T275[5];
  assign T905[4] = T282[4] | T275[4];
  assign T905[3] = T282[3] | T275[3];
  assign T905[2] = T282[2] | T275[2];
  assign T905[1] = T282[1] | T275[1];
  assign T905[0] = T282[0] | T275[0];
  assign N140 = ~T281;
  assign T280 = N327 | N330;
  assign T281 = cyc_A3_sqrt | N320;
  assign cyc_A3_sqrt = N330 & sqrtOp_PA;
  assign T282[20] = T295[20] | T283[20];
  assign T282[19] = T295[19] | T283[19];
  assign T282[18] = T295[18] | T283[18];
  assign T282[17] = T295[17] | T283[17];
  assign T282[16] = T295[16] | T283[16];
  assign T282[15] = T295[15] | T283[15];
  assign T282[14] = T295[14] | T283[14];
  assign T282[13] = T295[13] | T283[13];
  assign T282[12] = T295[12] | T283[12];
  assign T282[11] = T295[11] | T283[11];
  assign T282[10] = T295[10] | T283[10];
  assign T282[9] = T295[9] | T283[9];
  assign T282[8] = T295[8] | T283[8];
  assign T282[7] = T295[7] | T283[7];
  assign T282[6] = T295[6] | T283[6];
  assign T282[5] = T295[5] | T283[5];
  assign T282[4] = T295[4] | T283[4];
  assign T282[3] = T295[3] | T283[3];
  assign T282[2] = T295[2] | T283[2];
  assign T282[1] = T295[1] | T283[1];
  assign T282[0] = T295[0] | T283[0];
  assign N141 = ~T287;
  assign T287 = T289 | cyc_A3_div;
  assign cyc_A3_div = N330 & T288;
  assign T288 = ~sqrtOp_PA;
  assign T289 = N327 & T908[9];
  assign T295[20] = T300[20] | 1'b0;
  assign T295[19] = T300[19] | 1'b0;
  assign T295[18] = T300[18] | 1'b0;
  assign T295[17] = T300[17] | 1'b0;
  assign T295[16] = T300[16] | 1'b0;
  assign T295[15] = T300[15] | 1'b0;
  assign T295[14] = T300[14] | 1'b0;
  assign T295[13] = T300[13] | 1'b0;
  assign T295[12] = T300[12] | 1'b0;
  assign T295[11] = T300[11] | 1'b0;
  assign T295[10] = T300[10] | T910[10];
  assign T295[9] = T300[9] | 1'b0;
  assign T295[8] = T300[8] | 1'b0;
  assign T295[7] = T300[7] | 1'b0;
  assign T295[6] = T300[6] | 1'b0;
  assign T295[5] = T300[5] | 1'b0;
  assign T295[4] = T300[4] | 1'b0;
  assign T295[3] = T300[3] | 1'b0;
  assign T295[2] = T300[2] | 1'b0;
  assign T295[1] = T300[1] | 1'b0;
  assign T295[0] = T300[0] | 1'b0;
  assign T910[10] = T297;
  assign T297 = N327 & T298;
  assign T298 = ~T908[9];
  assign T300[20] = T304[20] | 1'b0;
  assign T300[19] = T304[19] | T911[19];
  assign T300[18] = T304[18] | T911[18];
  assign T300[17] = T304[17] | T911[17];
  assign T300[16] = T304[16] | T911[16];
  assign T300[15] = T304[15] | T911[15];
  assign T300[14] = T304[14] | T911[14];
  assign T300[13] = T304[13] | T911[13];
  assign T300[12] = T304[12] | T911[12];
  assign T300[11] = T304[11] | T911[11];
  assign T300[10] = T304[10] | T911[10];
  assign T300[9] = T304[9] | T911[9];
  assign T300[8] = T304[8] | T911[8];
  assign T300[7] = T304[7] | T911[7];
  assign T300[6] = T304[6] | T911[6];
  assign T300[5] = T304[5] | T911[5];
  assign T300[4] = T304[4] | T911[4];
  assign T300[3] = T304[3] | T911[3];
  assign T300[2] = T304[2] | T911[2];
  assign T300[1] = T304[1] | T911[1];
  assign T300[0] = T304[0] | T911[0];
  assign T304[20] = 1'b0 | T305[20];
  assign T304[19] = T914[19] | T305[19];
  assign T304[18] = T914[18] | T305[18];
  assign T304[17] = T914[17] | T305[17];
  assign T304[16] = T914[16] | T305[16];
  assign T304[15] = T914[15] | T305[15];
  assign T304[14] = T914[14] | T305[14];
  assign T304[13] = T914[13] | T305[13];
  assign T304[12] = T914[12] | T305[12];
  assign T304[11] = T914[11] | T305[11];
  assign T304[10] = T914[10] | T305[10];
  assign T304[9] = T914[9] | T305[9];
  assign T304[8] = T914[8] | T305[8];
  assign T304[7] = T914[7] | T305[7];
  assign T304[6] = T914[6] | T305[7];
  assign T304[5] = T914[5] | T305[7];
  assign T304[4] = T914[4] | T305[7];
  assign T304[3] = T914[3] | T305[7];
  assign T304[2] = T914[2] | T305[7];
  assign T304[1] = T914[1] | T305[7];
  assign T304[0] = T914[0] | T305_0;
  assign T305[19] = T311[11] | T308[11];
  assign T305[18] = T311[10] | T308[11];
  assign T305[17] = T311[9] | T308[11];
  assign T305[16] = T311[8] | 1'b0;
  assign T305[15] = T311[7] | T308[11];
  assign T305[14] = T311[6] | T308[11];
  assign T305[13] = T311[5] | T308[11];
  assign T305[12] = T311[4] | T308[11];
  assign T305[11] = T311[3] | 1'b0;
  assign T305[10] = T311[2] | T308[11];
  assign T305[9] = T311[1] | 1'b0;
  assign T305[8] = T311[0] | 1'b0;
  assign T308[11] = zLinPiece_7_A4_div;
  assign zLinPiece_7_A4_div = T305[20] & N332;
  assign T311[11] = T315[11] | T312[11];
  assign T311[10] = T315[10] | T312[11];
  assign T311[9] = T315[9] | 1'b0;
  assign T311[8] = T315[8] | T312[11];
  assign T311[7] = T315[7] | T312[11];
  assign T311[6] = T315[6] | 1'b0;
  assign T311[5] = T315[5] | T312[11];
  assign T311[4] = T315[4] | T312[11];
  assign T311[3] = T315[3] | T312[11];
  assign T311[2] = T315[2] | T312[11];
  assign T311[1] = T315[1] | 1'b0;
  assign T311[0] = T315[0] | T312[11];
  assign T312[11] = zLinPiece_6_A4_div;
  assign zLinPiece_6_A4_div = T305[20] & N337;
  assign T315[11] = T319[11] | T316[11];
  assign T315[10] = T319[10] | T316[11];
  assign T315[9] = T319[9] | 1'b0;
  assign T315[8] = T319[8] | 1'b0;
  assign T315[7] = T319[7] | 1'b0;
  assign T315[6] = T319[6] | T316[11];
  assign T315[5] = T319[5] | 1'b0;
  assign T315[4] = T319[4] | T316[11];
  assign T315[3] = T319[3] | 1'b0;
  assign T315[2] = T319[2] | T316[11];
  assign T315[1] = T319[1] | T316[11];
  assign T315[0] = T319[0] | 1'b0;
  assign T316[11] = zLinPiece_5_A4_div;
  assign zLinPiece_5_A4_div = T305[20] & N341;
  assign T319[11] = T323[11] | T320[11];
  assign T319[10] = T323[10] | 1'b0;
  assign T319[9] = T323[9] | T320[11];
  assign T319[8] = T323[8] | 1'b0;
  assign T319[7] = T323[7] | T320[11];
  assign T319[6] = T323[6] | 1'b0;
  assign T319[5] = T323[5] | T320[11];
  assign T319[4] = T323[4] | T320[11];
  assign T319[3] = T323[3] | 1'b0;
  assign T319[2] = T323[2] | T320[11];
  assign T319[1] = T323[1] | 1'b0;
  assign T319[0] = T323[0] | 1'b0;
  assign T320[11] = zLinPiece_4_A4_div;
  assign zLinPiece_4_A4_div = T305[20] & N343;
  assign T323[11] = T327[11] | T324[11];
  assign T323[10] = T327[10] | 1'b0;
  assign T323[9] = T327[9] | 1'b0;
  assign T323[8] = T327[8] | 1'b0;
  assign T323[7] = T327[7] | T324[11];
  assign T323[6] = T327[6] | T324[11];
  assign T323[5] = T327[5] | 1'b0;
  assign T323[4] = T327[4] | 1'b0;
  assign T323[3] = T327[3] | 1'b0;
  assign T323[2] = T327[2] | T324[11];
  assign T323[1] = T327[1] | T324[11];
  assign T323[0] = T327[0] | 1'b0;
  assign T324[11] = zLinPiece_3_A4_div;
  assign zLinPiece_3_A4_div = T305[20] & N346;
  assign T327[11] = T331[11] | 1'b0;
  assign T327[10] = T331[10] | T328[10];
  assign T327[9] = T331[9] | T328[10];
  assign T327[8] = T331[8] | 1'b0;
  assign T327[7] = T331[7] | 1'b0;
  assign T327[6] = T331[6] | T328[10];
  assign T327[5] = T331[5] | T328[10];
  assign T327[4] = T331[4] | T328[10];
  assign T327[3] = T331[3] | 1'b0;
  assign T327[2] = T331[2] | T328[10];
  assign T327[1] = T331[1] | 1'b0;
  assign T327[0] = T331[0] | T328[10];
  assign T328[10] = zLinPiece_2_A4_div;
  assign zLinPiece_2_A4_div = T305[20] & N351;
  assign T331[11] = 1'b0 | 1'b0;
  assign T331[10] = 1'b0 | 1'b0;
  assign T331[9] = 1'b0 | T332[9];
  assign T331[8] = 1'b0 | T332[9];
  assign T331[7] = 1'b0 | T332[9];
  assign T331[6] = 1'b0 | 1'b0;
  assign T331[5] = 1'b0 | T332[9];
  assign T331[4] = T335[4] | 1'b0;
  assign T331[3] = T335[4] | 1'b0;
  assign T331[2] = T335[4] | 1'b0;
  assign T331[1] = 1'b0 | T332[9];
  assign T331[0] = 1'b0 | 1'b0;
  assign T332[9] = zLinPiece_1_A4_div;
  assign zLinPiece_1_A4_div = T305[20] & N356;
  assign T335[4] = zLinPiece_0_A4_div;
  assign zLinPiece_0_A4_div = T305[20] & N354;
  assign T914[19] = T364[19] | N349;
  assign T914[18] = T364[18] | T339[18];
  assign T914[17] = T364[17] | T339[17];
  assign T914[16] = T364[16] | T339[16];
  assign T914[15] = T364[15] | T339[15];
  assign T914[14] = T364[14] | T339[14];
  assign T914[13] = T364[13] | T339[13];
  assign T914[12] = T364[12] | T339[12];
  assign T914[11] = T364[11] | T339[11];
  assign T914[10] = T364[10] | T339[10];
  assign T914[9] = 1'b0 | T339[9];
  assign T914[8] = 1'b0 | T339[8];
  assign T914[7] = 1'b0 | T339[7];
  assign T914[6] = 1'b0 | T339[6];
  assign T914[5] = 1'b0 | T339[5];
  assign T914[4] = 1'b0 | T339[5];
  assign T914[3] = 1'b0 | T339[5];
  assign T914[2] = 1'b0 | T339[5];
  assign T914[1] = 1'b0 | T339[5];
  assign T914[0] = 1'b0 | T339_0;
  assign T339[18] = T346[12] | T342[12];
  assign T339[17] = T346[11] | T342[12];
  assign T339[16] = T346[10] | 1'b0;
  assign T339[15] = T346[9] | T342[12];
  assign T339[14] = T346[8] | T342[12];
  assign T339[13] = T346[7] | 1'b0;
  assign T339[12] = T346[6] | 1'b0;
  assign T339[11] = T346[5] | 1'b0;
  assign T339[10] = T346[4] | T342[12];
  assign T339[9] = T346[3] | 1'b0;
  assign T339[8] = T346[2] | T342[12];
  assign T339[7] = T346[1] | T342[12];
  assign T339[6] = T346[0] | T342[12];
  assign T342[12] = zQuadPiece_3_A6_sqrt;
  assign zQuadPiece_3_A6_sqrt = T344 & sigB_PA_51;
  assign T344 = N349 & exp_PA[0];
  assign T346[12] = T352[12] | T347[12];
  assign T346[11] = T352[11] | 1'b0;
  assign T346[10] = T352[10] | 1'b0;
  assign T346[9] = T352[9] | T347[12];
  assign T346[8] = T352[8] | 1'b0;
  assign T346[7] = T352[7] | T347[12];
  assign T346[6] = T352[6] | T347[12];
  assign T346[5] = T352[5] | 1'b0;
  assign T346[4] = T352[4] | T347[12];
  assign T346[3] = T352[3] | 1'b0;
  assign T346[2] = T352[2] | 1'b0;
  assign T346[1] = T352[1] | T347[12];
  assign T346[0] = T352[0] | T347[12];
  assign T347[12] = zQuadPiece_2_A6_sqrt;
  assign zQuadPiece_2_A6_sqrt = T350 & T348;
  assign T348 = ~sigB_PA_51;
  assign T350 = N349 & exp_PA[0];
  assign T352[12] = 1'b0 | 1'b0;
  assign T352[11] = 1'b0 | T353[11];
  assign T352[10] = 1'b0 | 1'b0;
  assign T352[9] = 1'b0 | T353[11];
  assign T352[8] = 1'b0 | T353[11];
  assign T352[7] = 1'b0 | T353[11];
  assign T352[6] = 1'b0 | T353[11];
  assign T352[5] = 1'b0 | 1'b0;
  assign T352[4] = T358[4] | 1'b0;
  assign T352[3] = T358[4] | T353[11];
  assign T352[2] = 1'b0 | 1'b0;
  assign T352[1] = T358[4] | T353[11];
  assign T352[0] = 1'b0 | 1'b0;
  assign T353[11] = zQuadPiece_1_A6_sqrt;
  assign zQuadPiece_1_A6_sqrt = T355 & sigB_PA_51;
  assign T355 = N349 & T356;
  assign T356 = ~exp_PA[0];
  assign T358[4] = zQuadPiece_0_A6_sqrt;
  assign zQuadPiece_0_A6_sqrt = T361 & T359;
  assign T359 = ~sigB_PA_51;
  assign T361 = N349 & T362;
  assign T362 = ~exp_PA[0];
  assign T364[19] = T369[9] | T365[9];
  assign T364[18] = T369[8] | 1'b0;
  assign T364[17] = T369[7] | 1'b0;
  assign T364[16] = T369[6] | T365[9];
  assign T364[15] = T369[5] | T365[9];
  assign T364[14] = T369[4] | T365[9];
  assign T364[13] = T369[3] | T365[9];
  assign T364[12] = T369[2] | T365[9];
  assign T364[11] = T369[1] | T365[9];
  assign T364[10] = T369[0] | 1'b0;
  assign T365[9] = zQuadPiece_3_A7_sqrt;
  assign zQuadPiece_3_A7_sqrt = T367 & io_b[51];
  assign T367 = cyc_A7_sqrt & io_b[52];
  assign T369[9] = T375[9] | 1'b0;
  assign T369[8] = T375[8] | T370[8];
  assign T369[7] = T375[7] | 1'b0;
  assign T369[6] = T375[6] | T370[8];
  assign T369[5] = T375[5] | 1'b0;
  assign T369[4] = T375[4] | 1'b0;
  assign T369[3] = T375[3] | T370[8];
  assign T369[2] = T375[2] | T370[8];
  assign T369[1] = T375[1] | 1'b0;
  assign T369[0] = T375[0] | T370[8];
  assign T370[8] = zQuadPiece_2_A7_sqrt;
  assign zQuadPiece_2_A7_sqrt = T373 & T371;
  assign T371 = ~io_b[51];
  assign T373 = cyc_A7_sqrt & io_b[52];
  assign T375[9] = 1'b0 | 1'b0;
  assign T375[8] = 1'b0 | T376[8];
  assign T375[7] = 1'b0 | T376[8];
  assign T375[6] = 1'b0 | T376[8];
  assign T375[5] = T381[5] | 1'b0;
  assign T375[4] = 1'b0 | T376[8];
  assign T375[3] = T381[5] | T376[8];
  assign T375[2] = T381[5] | T376[8];
  assign T375[1] = T381[5] | T376[8];
  assign T375[0] = T381[5] | T376[8];
  assign T376[8] = zQuadPiece_1_A7_sqrt;
  assign zQuadPiece_1_A7_sqrt = T378 & io_b[51];
  assign T378 = cyc_A7_sqrt & T379;
  assign T379 = ~io_b[52];
  assign T381[5] = zQuadPiece_0_A7_sqrt;
  assign zQuadPiece_0_A7_sqrt = T384 & T382;
  assign T382 = ~io_b[51];
  assign T384 = cyc_A7_sqrt & T385;
  assign T385 = ~io_b[52];
  assign mulAdd9B_A[8] = T408[8] | T388[8];
  assign mulAdd9B_A[7] = T408[7] | T388[7];
  assign mulAdd9B_A[6] = T408[6] | T388[6];
  assign mulAdd9B_A[5] = T408[5] | T388[5];
  assign mulAdd9B_A[4] = T408[4] | T388[4];
  assign mulAdd9B_A[3] = T408[3] | T388[3];
  assign mulAdd9B_A[2] = T408[2] | T388[2];
  assign mulAdd9B_A[1] = T408[1] | T388[1];
  assign mulAdd9B_A[0] = T408[0] | T388[0];
  assign N142 = ~T407;
  assign T390[8] = T394[8] | T391[8];
  assign T390[7] = T394[7] | T391[7];
  assign T390[6] = T394[6] | T391[6];
  assign T390[5] = T394[5] | T391[5];
  assign T390[4] = T394[4] | T391[4];
  assign T390[3] = T394[3] | T391[3];
  assign T390[2] = T394[2] | T391[2];
  assign T390[1] = T394[1] | T391[1];
  assign T390[0] = T394[0] | T391[0];
  assign T391[8] = N320;
  assign T394[8] = T397[8] | T395[8];
  assign T394[7] = T397[7] | T395[7];
  assign T394[6] = T397[6] | T395[6];
  assign T394[5] = T397[5] | T395[5];
  assign T394[4] = T397[4] | T395[4];
  assign T394[3] = T397[3] | T395[3];
  assign T394[2] = T397[2] | T395[2];
  assign T394[1] = T397[1] | T395[1];
  assign T394[0] = T397[0] | T395[0];
  assign T397[8] = T398[8] | zFractR0_A4_div[8];
  assign T397[7] = T398[7] | zFractR0_A4_div[7];
  assign T397[6] = T398[6] | zFractR0_A4_div[6];
  assign T397[5] = T398[5] | zFractR0_A4_div[5];
  assign T397[4] = T398[4] | zFractR0_A4_div[4];
  assign T397[3] = T398[3] | zFractR0_A4_div[3];
  assign T397[2] = T398[2] | zFractR0_A4_div[2];
  assign T397[1] = T398[1] | zFractR0_A4_div[1];
  assign T397[0] = T398[0] | zFractR0_A4_div[0];
  assign T398[8] = T401[8] | T399[8];
  assign T398[7] = T401[7] | T399[7];
  assign T398[6] = T401[6] | T399[6];
  assign T398[5] = T401[5] | T399[5];
  assign T398[4] = T401[4] | T399[4];
  assign T398[3] = T401[3] | T399[3];
  assign T398[2] = T401[2] | T399[2];
  assign T398[1] = T401[1] | T399[1];
  assign T398[0] = T401[0] | T399[0];
  assign T401[8] = T402[8] | zFractR0_A6_sqrt[8];
  assign T401[7] = T402[7] | zFractR0_A6_sqrt[7];
  assign T401[6] = T402[6] | zFractR0_A6_sqrt[6];
  assign T401[5] = T402[5] | zFractR0_A6_sqrt[5];
  assign T401[4] = T402[4] | zFractR0_A6_sqrt[4];
  assign T401[3] = T402[3] | zFractR0_A6_sqrt[3];
  assign T401[2] = T402[2] | zFractR0_A6_sqrt[2];
  assign T401[1] = T402[1] | zFractR0_A6_sqrt[1];
  assign T401[0] = T402[0] | zFractR0_A6_sqrt[0];
  assign N143 = ~cyc_A7_sqrt;
  assign T403 = T404 | N320;
  assign T404 = T405 | cyc_A4;
  assign cyc_A4 = N327 | T305[20];
  assign T405 = T406 | N324;
  assign T406 = cyc_A7_sqrt | N349;
  assign T407 = ~cyc_S;
  assign T408[8] = zK1_A4_div[8] | T402[8];
  assign T408[7] = zK1_A4_div[7] | T402[7];
  assign T408[6] = zK1_A4_div[6] | T402[6];
  assign T408[5] = zK1_A4_div[5] | T402[5];
  assign T408[4] = zK1_A4_div[4] | T402[4];
  assign T408[3] = zK1_A4_div[3] | T402[3];
  assign T408[2] = zK1_A4_div[2] | T402[2];
  assign T408[1] = zK1_A4_div[1] | T402[1];
  assign T408[0] = zK1_A4_div[0] | T402[0];
  assign zK1_A4_div[8] = T411[8] | 1'b0;
  assign zK1_A4_div[7] = T411[7] | T410[7];
  assign zK1_A4_div[6] = T411[6] | 1'b0;
  assign zK1_A4_div[5] = T411[5] | 1'b0;
  assign zK1_A4_div[4] = T411[4] | 1'b0;
  assign zK1_A4_div[3] = T411[3] | T410[7];
  assign zK1_A4_div[2] = T411[2] | 1'b0;
  assign zK1_A4_div[1] = T411[1] | 1'b0;
  assign zK1_A4_div[0] = T411[0] | T410[7];
  assign T410[7] = zLinPiece_7_A4_div;
  assign T411[8] = T413[8] | 1'b0;
  assign T411[7] = T413[7] | T412[7];
  assign T411[6] = T413[6] | 1'b0;
  assign T411[5] = T413[5] | 1'b0;
  assign T411[4] = T413[4] | T412[7];
  assign T411[3] = T413[3] | T412[7];
  assign T411[2] = T413[2] | T412[7];
  assign T411[1] = T413[1] | 1'b0;
  assign T411[0] = T413[0] | 1'b0;
  assign T412[7] = zLinPiece_6_A4_div;
  assign T413[8] = T415[8] | 1'b0;
  assign T413[7] = T415[7] | T414[7];
  assign T413[6] = T415[6] | 1'b0;
  assign T413[5] = T415[5] | T414[7];
  assign T413[4] = T415[4] | T414[7];
  assign T413[3] = T415[3] | 1'b0;
  assign T413[2] = T415[2] | T414[7];
  assign T413[1] = T415[1] | 1'b0;
  assign T413[0] = T415[0] | 1'b0;
  assign T414[7] = zLinPiece_5_A4_div;
  assign T415[8] = T417[8] | 1'b0;
  assign T415[7] = T417[7] | T416[7];
  assign T415[6] = T417[6] | T416[7];
  assign T415[5] = T417[5] | 1'b0;
  assign T415[4] = T417[4] | T416[7];
  assign T415[3] = T417[3] | 1'b0;
  assign T415[2] = T417[2] | 1'b0;
  assign T415[1] = T417[1] | T416[7];
  assign T415[0] = T417[0] | 1'b0;
  assign T416[7] = zLinPiece_4_A4_div;
  assign T417[8] = T419[8] | 1'b0;
  assign T417[7] = T419[7] | T418[7];
  assign T417[6] = T419[6] | T418[7];
  assign T417[5] = T419[5] | T418[7];
  assign T417[4] = T419[4] | T418[7];
  assign T417[3] = T419[3] | T418[7];
  assign T417[2] = T419[2] | 1'b0;
  assign T417[1] = T419[1] | 1'b0;
  assign T417[0] = T419[0] | 1'b0;
  assign T418[7] = zLinPiece_3_A4_div;
  assign T419[8] = T421[8] | T420[8];
  assign T419[7] = T421[7] | 1'b0;
  assign T419[6] = T421[6] | 1'b0;
  assign T419[5] = T421[5] | T420[8];
  assign T419[4] = T421[4] | 1'b0;
  assign T419[3] = T421[3] | T420[8];
  assign T419[2] = T421[2] | 1'b0;
  assign T419[1] = T421[1] | T420[8];
  assign T419[0] = T421[0] | 1'b0;
  assign T420[8] = zLinPiece_2_A4_div;
  assign T421[8] = T423[8] | T422[8];
  assign T421[7] = T423[8] | 1'b0;
  assign T421[6] = T423[8] | T422[8];
  assign T421[5] = 1'b0 | T422[8];
  assign T421[4] = 1'b0 | 1'b0;
  assign T421[3] = 1'b0 | T422[8];
  assign T421[2] = T423[8] | T422[8];
  assign T421[1] = T423[8] | 1'b0;
  assign T421[0] = T423[8] | 1'b0;
  assign T422[8] = zLinPiece_1_A4_div;
  assign T423[8] = zLinPiece_0_A4_div;
  assign mulAdd9A_A[8] = T451[8] | T424[8];
  assign mulAdd9A_A[7] = T451[7] | T424[7];
  assign mulAdd9A_A[6] = T451[6] | T424[6];
  assign mulAdd9A_A[5] = T451[5] | T424[5];
  assign mulAdd9A_A[4] = T451[4] | T424[4];
  assign mulAdd9A_A[3] = T451[3] | T424[3];
  assign mulAdd9A_A[2] = T451[2] | T424[2];
  assign mulAdd9A_A[1] = T451[1] | T424[1];
  assign mulAdd9A_A[0] = T451[0] | T424[0];
  assign N144 = ~T450;
  assign N145 = ~T445;
  assign T426[8] = T432[8] | T919[8];
  assign T426[7] = T432[7] | T919[7];
  assign T426[6] = T432[6] | T919[6];
  assign T426[5] = T432[5] | T919[5];
  assign T426[4] = T432[4] | T919[4];
  assign T426[3] = T432[3] | T919[3];
  assign T426[2] = T432[2] | T919[2];
  assign T426[1] = T432[1] | T919[1];
  assign T426[0] = T432[0] | T919[0];
  assign N146 = ~T430;
  assign T428[8] = ~T251[1];
  assign T428[7] = ~T251[0];
  assign T428[6] = ~mulAdd9Out_A[8];
  assign T428[5] = ~mulAdd9Out_A[7];
  assign T428[4] = ~mulAdd9Out_A[6];
  assign T428[3] = ~mulAdd9Out_A[5];
  assign T428[2] = ~mulAdd9Out_A[4];
  assign T428[1] = ~mulAdd9Out_A[3];
  assign T428[0] = ~mulAdd9Out_A[2];
  assign T430 = N320 & T251[2];
  assign T432[8] = T436[8] | T920[8];
  assign T432[7] = T436[7] | T920[7];
  assign T432[6] = T436[6] | T920[6];
  assign T432[5] = T436[5] | T920[5];
  assign T432[4] = T436[4] | T920[4];
  assign T432[3] = T436[3] | T920[3];
  assign T432[2] = T436[2] | T920[2];
  assign T432[1] = T436[1] | T920[1];
  assign T432[0] = T436[0] | T920[0];
  assign N147 = ~T435;
  assign T920[8] = T435;
  assign T435 = N324 | N330;
  assign T436[8] = T438[8] | T921[8];
  assign T436[7] = T438[7] | T921[7];
  assign T436[6] = T438[6] | T921[6];
  assign T436[5] = T438[5] | T921[5];
  assign T436[4] = T438[4] | T921[4];
  assign T436[3] = T438[3] | T921[3];
  assign T436[2] = T438[2] | T921[2];
  assign T436[1] = T438[1] | T921[1];
  assign T436[0] = T438[0] | T921[0];
  assign N148 = ~T305[20];
  assign T438[8] = T441[8] | T922[8];
  assign T438[7] = T441[7] | T922[7];
  assign T438[6] = T441[6] | T922[6];
  assign T438[5] = T441[5] | T922[5];
  assign T438[4] = T441[4] | T922[4];
  assign T438[3] = T441[3] | T922[3];
  assign T438[2] = T441[2] | T922[2];
  assign T438[1] = T441[1] | T922[1];
  assign T438[0] = T441[0] | T922[0];
  assign T441[8] = T442[8] | zFractR0_A6_sqrt[8];
  assign T441[7] = T442[7] | zFractR0_A6_sqrt[7];
  assign T441[6] = T442[6] | zFractR0_A6_sqrt[6];
  assign T441[5] = T442[5] | zFractR0_A6_sqrt[5];
  assign T441[4] = T442[4] | zFractR0_A6_sqrt[4];
  assign T441[3] = T442[3] | zFractR0_A6_sqrt[3];
  assign T441[2] = T442[2] | zFractR0_A6_sqrt[2];
  assign T441[1] = T442[1] | zFractR0_A6_sqrt[1];
  assign T441[0] = T442[0] | zFractR0_A6_sqrt[0];
  assign T443[8] = ~T251[10];
  assign T443[7] = ~T251[9];
  assign T443[6] = ~T251[8];
  assign T443[5] = ~T251[7];
  assign T443[4] = ~T251[6];
  assign T443[3] = ~T251[5];
  assign T443[2] = ~T251[4];
  assign T443[1] = ~T251[3];
  assign T443[0] = ~T251[2];
  assign T445 = T446 | N320;
  assign T446 = T447 | N330;
  assign T447 = T448 | cyc_A4;
  assign T448 = T449 | N324;
  assign T449 = cyc_A7_sqrt | N349;
  assign T450 = ~cyc_S;
  assign T451[8] = zFractB_A4_div[48] | zK2_A7_sqrt[8];
  assign T451[7] = zFractB_A4_div[47] | zK2_A7_sqrt[7];
  assign T451[6] = zFractB_A4_div[46] | zK2_A7_sqrt[6];
  assign T451[5] = zFractB_A4_div[45] | zK2_A7_sqrt[5];
  assign T451[4] = zFractB_A4_div[44] | zK2_A7_sqrt[4];
  assign T451[3] = T921[8] | zK2_A7_sqrt[3];
  assign T451[2] = T921[7] | zK2_A7_sqrt[2];
  assign T451[1] = T921[6] | zK2_A7_sqrt[1];
  assign T451[0] = T921[5] | zK2_A7_sqrt[0];
  assign zK2_A7_sqrt[8] = T453[8] | 1'b0;
  assign zK2_A7_sqrt[7] = T453[7] | T452[7];
  assign zK2_A7_sqrt[6] = T453[6] | 1'b0;
  assign zK2_A7_sqrt[5] = T453[5] | 1'b0;
  assign zK2_A7_sqrt[4] = T453[4] | 1'b0;
  assign zK2_A7_sqrt[3] = T453[3] | T452[7];
  assign zK2_A7_sqrt[2] = T453[2] | 1'b0;
  assign zK2_A7_sqrt[1] = T453[1] | 1'b0;
  assign zK2_A7_sqrt[0] = T453[0] | T452[7];
  assign T452[7] = zQuadPiece_3_A7_sqrt;
  assign T453[8] = T455[8] | T454[8];
  assign T453[7] = T455[7] | 1'b0;
  assign T453[6] = T455[6] | T454[8];
  assign T453[5] = T455[5] | 1'b0;
  assign T453[4] = T455[4] | 1'b0;
  assign T453[3] = T455[3] | 1'b0;
  assign T453[2] = T455[2] | 1'b0;
  assign T453[1] = T455[1] | T454[8];
  assign T453[0] = T455[0] | T454[8];
  assign T454[8] = zQuadPiece_2_A7_sqrt;
  assign T455[8] = T457[8] | 1'b0;
  assign T455[7] = T457[8] | T456[7];
  assign T455[6] = T457[8] | T456[7];
  assign T455[5] = 1'b0 | 1'b0;
  assign T455[4] = 1'b0 | 1'b0;
  assign T455[3] = T457[8] | 1'b0;
  assign T455[2] = 1'b0 | 1'b0;
  assign T455[1] = 1'b0 | 1'b0;
  assign T455[0] = 1'b0 | T456[7];
  assign T456[7] = zQuadPiece_1_A7_sqrt;
  assign T457[8] = zQuadPiece_0_A7_sqrt;
  assign N149 = ~loMulAdd9Out_A[18];
  assign cyc_A1_sqrt = N316 & sqrtOp_PA;
  assign cyc_B6_sqrt = T468 & sqrtOp_PB;
  assign T468 = N502 & valid_PB;
  assign T925[51] = T475[51] | 1'b0;
  assign T925[50] = T475[50] | T926[50];
  assign T925[49] = T475[49] | T926[49];
  assign T925[48] = T475[48] | T926[48];
  assign T925[47] = T475[47] | T926[47];
  assign T925[46] = T475[46] | T926[46];
  assign T925[45] = T475[45] | T926[45];
  assign T925[44] = T475[44] | T926[44];
  assign T925[43] = T475[43] | T926[43];
  assign T925[42] = T475[42] | T926[42];
  assign T925[41] = T475[41] | T926[41];
  assign T925[40] = T475[40] | T926[40];
  assign T925[39] = T475[39] | T926[39];
  assign T925[38] = T475[38] | T926[38];
  assign T925[37] = T475[37] | T926[37];
  assign T925[36] = T475[36] | T926[36];
  assign T925[35] = 1'b0 | T926[35];
  assign T925[34] = 1'b0 | T926[34];
  assign T925[33] = 1'b0 | T926[33];
  assign T925[32] = 1'b0 | T926[32];
  assign T925[31] = 1'b0 | T926[31];
  assign T925[30] = 1'b0 | T926[30];
  assign T925[29] = 1'b0 | T926[29];
  assign T925[28] = 1'b0 | T926[28];
  assign T925[27] = 1'b0 | T926[27];
  assign T925[26] = 1'b0 | T926[26];
  assign T925[25] = 1'b0 | T926[25];
  assign T925[24] = 1'b0 | T926[24];
  assign T925[23] = 1'b0 | T926[23];
  assign T925[22] = 1'b0 | T926[22];
  assign T925[21] = 1'b0 | T926[21];
  assign T925[20] = 1'b0 | T926[20];
  assign T925[19] = 1'b0 | T926[19];
  assign T925[18] = 1'b0 | 1'b0;
  assign T925[17] = 1'b0 | 1'b0;
  assign T925[16] = 1'b0 | 1'b0;
  assign T925[15] = 1'b0 | 1'b0;
  assign T925[14] = 1'b0 | 1'b0;
  assign T925[13] = 1'b0 | 1'b0;
  assign T925[12] = 1'b0 | 1'b0;
  assign T925[11] = 1'b0 | 1'b0;
  assign T925[10] = 1'b0 | 1'b0;
  assign T925[9] = 1'b0 | 1'b0;
  assign T925[8] = 1'b0 | 1'b0;
  assign T925[7] = 1'b0 | 1'b0;
  assign T925[6] = 1'b0 | 1'b0;
  assign T925[5] = 1'b0 | 1'b0;
  assign T925[4] = 1'b0 | 1'b0;
  assign T925[3] = 1'b0 | 1'b0;
  assign T925[2] = 1'b0 | 1'b0;
  assign T925[1] = 1'b0 | 1'b0;
  assign T925[0] = 1'b0 | 1'b0;
  assign io_latchMulAddB_0 = T478 | N312;
  assign T478 = T479 | N476;
  assign T479 = T480 | N308;
  assign T480 = T481 | N513;
  assign T481 = T482 | cyc_B6_sqrt;
  assign T482 = N316 | N506;
  assign io_mulAddA_0[53] = 1'b0 | zComplSigT_C1_sqrt[53];
  assign io_mulAddA_0[52] = T927[52] | zComplSigT_C1_sqrt[52];
  assign io_mulAddA_0[51] = T927[51] | zComplSigT_C1_sqrt[51];
  assign io_mulAddA_0[50] = T927[50] | zComplSigT_C1_sqrt[50];
  assign io_mulAddA_0[49] = T927[49] | zComplSigT_C1_sqrt[49];
  assign io_mulAddA_0[48] = T927[48] | zComplSigT_C1_sqrt[48];
  assign io_mulAddA_0[47] = T927[47] | zComplSigT_C1_sqrt[47];
  assign io_mulAddA_0[46] = T927[46] | zComplSigT_C1_sqrt[46];
  assign io_mulAddA_0[45] = T927[45] | zComplSigT_C1_sqrt[45];
  assign io_mulAddA_0[44] = T927[44] | zComplSigT_C1_sqrt[44];
  assign io_mulAddA_0[43] = T927[43] | zComplSigT_C1_sqrt[43];
  assign io_mulAddA_0[42] = T927[42] | zComplSigT_C1_sqrt[42];
  assign io_mulAddA_0[41] = T927[41] | zComplSigT_C1_sqrt[41];
  assign io_mulAddA_0[40] = T927[40] | zComplSigT_C1_sqrt[40];
  assign io_mulAddA_0[39] = T927[39] | zComplSigT_C1_sqrt[39];
  assign io_mulAddA_0[38] = T927[38] | zComplSigT_C1_sqrt[38];
  assign io_mulAddA_0[37] = T927[37] | zComplSigT_C1_sqrt[37];
  assign io_mulAddA_0[36] = T927[36] | zComplSigT_C1_sqrt[36];
  assign io_mulAddA_0[35] = T927[35] | zComplSigT_C1_sqrt[35];
  assign io_mulAddA_0[34] = T927[34] | zComplSigT_C1_sqrt[34];
  assign io_mulAddA_0[33] = T927[33] | zComplSigT_C1_sqrt[33];
  assign io_mulAddA_0[32] = T927[32] | zComplSigT_C1_sqrt[32];
  assign io_mulAddA_0[31] = T927[31] | zComplSigT_C1_sqrt[31];
  assign io_mulAddA_0[30] = T927[30] | zComplSigT_C1_sqrt[30];
  assign io_mulAddA_0[29] = T927[29] | zComplSigT_C1_sqrt[29];
  assign io_mulAddA_0[28] = T927[28] | zComplSigT_C1_sqrt[28];
  assign io_mulAddA_0[27] = T927[27] | zComplSigT_C1_sqrt[27];
  assign io_mulAddA_0[26] = T927[26] | zComplSigT_C1_sqrt[26];
  assign io_mulAddA_0[25] = T927[25] | zComplSigT_C1_sqrt[25];
  assign io_mulAddA_0[24] = T927[24] | zComplSigT_C1_sqrt[24];
  assign io_mulAddA_0[23] = T927[23] | zComplSigT_C1_sqrt[23];
  assign io_mulAddA_0[22] = T927[22] | zComplSigT_C1_sqrt[22];
  assign io_mulAddA_0[21] = T927[21] | zComplSigT_C1_sqrt[21];
  assign io_mulAddA_0[20] = T927[20] | zComplSigT_C1_sqrt[20];
  assign io_mulAddA_0[19] = T927[19] | zComplSigT_C1_sqrt[19];
  assign io_mulAddA_0[18] = T927[18] | zComplSigT_C1_sqrt[18];
  assign io_mulAddA_0[17] = T927[17] | zComplSigT_C1_sqrt[17];
  assign io_mulAddA_0[16] = T927[16] | zComplSigT_C1_sqrt[16];
  assign io_mulAddA_0[15] = T927[15] | zComplSigT_C1_sqrt[15];
  assign io_mulAddA_0[14] = T927[14] | zComplSigT_C1_sqrt[14];
  assign io_mulAddA_0[13] = T927[13] | zComplSigT_C1_sqrt[13];
  assign io_mulAddA_0[12] = T927[12] | zComplSigT_C1_sqrt[12];
  assign io_mulAddA_0[11] = T927[11] | zComplSigT_C1_sqrt[11];
  assign io_mulAddA_0[10] = T927[10] | zComplSigT_C1_sqrt[10];
  assign io_mulAddA_0[9] = T927[9] | zComplSigT_C1_sqrt[9];
  assign io_mulAddA_0[8] = T927[8] | zComplSigT_C1_sqrt[8];
  assign io_mulAddA_0[7] = T927[7] | zComplSigT_C1_sqrt[7];
  assign io_mulAddA_0[6] = T927[6] | zComplSigT_C1_sqrt[6];
  assign io_mulAddA_0[5] = T927[5] | zComplSigT_C1_sqrt[5];
  assign io_mulAddA_0[4] = T927[4] | zComplSigT_C1_sqrt[4];
  assign io_mulAddA_0[3] = T927[3] | zComplSigT_C1_sqrt[3];
  assign io_mulAddA_0[2] = T927[2] | zComplSigT_C1_sqrt[2];
  assign io_mulAddA_0[1] = T927[1] | zComplSigT_C1_sqrt[1];
  assign io_mulAddA_0[0] = T927[0] | zComplSigT_C1_sqrt[0];
  assign N150 = ~cyc_C1_sqrt;
  assign T485[53] = ~io_mulAddResult_3[104];
  assign T485[52] = ~io_mulAddResult_3[103];
  assign T485[51] = ~io_mulAddResult_3[102];
  assign T485[50] = ~io_mulAddResult_3[101];
  assign T485[49] = ~io_mulAddResult_3[100];
  assign T485[48] = ~io_mulAddResult_3[99];
  assign T485[47] = ~io_mulAddResult_3[98];
  assign T485[46] = ~io_mulAddResult_3[97];
  assign T485[45] = ~io_mulAddResult_3[96];
  assign T485[44] = ~io_mulAddResult_3[95];
  assign T485[43] = ~io_mulAddResult_3[94];
  assign T485[42] = ~io_mulAddResult_3[93];
  assign T485[41] = ~io_mulAddResult_3[92];
  assign T485[40] = ~io_mulAddResult_3[91];
  assign T485[39] = ~io_mulAddResult_3[90];
  assign T485[38] = ~io_mulAddResult_3[89];
  assign T485[37] = ~io_mulAddResult_3[88];
  assign T485[36] = ~io_mulAddResult_3[87];
  assign T485[35] = ~io_mulAddResult_3[86];
  assign T485[34] = ~io_mulAddResult_3[85];
  assign T485[33] = ~io_mulAddResult_3[84];
  assign T485[32] = ~io_mulAddResult_3[83];
  assign T485[31] = ~io_mulAddResult_3[82];
  assign T485[30] = ~io_mulAddResult_3[81];
  assign T485[29] = ~io_mulAddResult_3[80];
  assign T485[28] = ~io_mulAddResult_3[79];
  assign T485[27] = ~io_mulAddResult_3[78];
  assign T485[26] = ~io_mulAddResult_3[77];
  assign T485[25] = ~io_mulAddResult_3[76];
  assign T485[24] = ~io_mulAddResult_3[75];
  assign T485[23] = ~io_mulAddResult_3[74];
  assign T485[22] = ~io_mulAddResult_3[73];
  assign T485[21] = ~io_mulAddResult_3[72];
  assign T485[20] = ~io_mulAddResult_3[71];
  assign T485[19] = ~io_mulAddResult_3[70];
  assign T485[18] = ~io_mulAddResult_3[69];
  assign T485[17] = ~io_mulAddResult_3[68];
  assign T485[16] = ~io_mulAddResult_3[67];
  assign T485[15] = ~io_mulAddResult_3[66];
  assign T485[14] = ~io_mulAddResult_3[65];
  assign T485[13] = ~io_mulAddResult_3[64];
  assign T485[12] = ~io_mulAddResult_3[63];
  assign T485[11] = ~io_mulAddResult_3[62];
  assign T485[10] = ~io_mulAddResult_3[61];
  assign T485[9] = ~io_mulAddResult_3[60];
  assign T485[8] = ~io_mulAddResult_3[59];
  assign T485[7] = ~io_mulAddResult_3[58];
  assign T485[6] = ~io_mulAddResult_3[57];
  assign T485[5] = ~io_mulAddResult_3[56];
  assign T485[4] = ~io_mulAddResult_3[55];
  assign T485[3] = ~io_mulAddResult_3[54];
  assign T485[2] = ~io_mulAddResult_3[53];
  assign T485[1] = ~io_mulAddResult_3[52];
  assign T485[0] = ~io_mulAddResult_3[51];
  assign T927[52] = T489[52] | T488[52];
  assign T927[51] = T489[51] | T488[51];
  assign T927[50] = T489[50] | T488[50];
  assign T927[49] = T489[49] | T488[49];
  assign T927[48] = T489[48] | T488[48];
  assign T927[47] = T489[47] | T488[47];
  assign T927[46] = T489[46] | T488[46];
  assign T927[45] = T489[45] | T488[45];
  assign T927[44] = T489[44] | T488[44];
  assign T927[43] = T489[43] | T488[43];
  assign T927[42] = T489[42] | T488[42];
  assign T927[41] = T489[41] | T488[41];
  assign T927[40] = T489[40] | T488[40];
  assign T927[39] = T489[39] | T488[39];
  assign T927[38] = T489[38] | T488[38];
  assign T927[37] = T489[37] | T488[37];
  assign T927[36] = T489[36] | T488[36];
  assign T927[35] = T489[35] | T488[35];
  assign T927[34] = T489[34] | T488[34];
  assign T927[33] = T489[33] | T488[33];
  assign T927[32] = T489[32] | T488[32];
  assign T927[31] = T489[31] | T488[31];
  assign T927[30] = T489[30] | T488[30];
  assign T927[29] = T489[29] | T488[29];
  assign T927[28] = T489[28] | T488[28];
  assign T927[27] = T489[27] | T488[27];
  assign T927[26] = T489[26] | T488[26];
  assign T927[25] = T489[25] | T488[25];
  assign T927[24] = T489[24] | T488[24];
  assign T927[23] = T489[23] | T488[23];
  assign T927[22] = T489[22] | T488[22];
  assign T927[21] = T489[21] | T488[21];
  assign T927[20] = T489[20] | T488[20];
  assign T927[19] = T489[19] | T488[19];
  assign T927[18] = T489[18] | T488[18];
  assign T927[17] = T489[17] | T488[17];
  assign T927[16] = T489[16] | T488[16];
  assign T927[15] = T489[15] | T488[15];
  assign T927[14] = T489[14] | T488[14];
  assign T927[13] = T489[13] | T488[13];
  assign T927[12] = T489[12] | T488[12];
  assign T927[11] = T489[11] | T488[11];
  assign T927[10] = T489[10] | T488[10];
  assign T927[9] = T489[9] | T488[9];
  assign T927[8] = T489[8] | T488[8];
  assign T927[7] = T489[7] | T488[7];
  assign T927[6] = T489[6] | T488[6];
  assign T927[5] = T489[5] | T488[5];
  assign T927[4] = T489[4] | T488[4];
  assign T927[3] = T489[3] | T488[3];
  assign T927[2] = T489[2] | T488[2];
  assign T927[1] = T489[1] | T488[1];
  assign T927[0] = T489[0] | T488[0];
  assign N151 = ~cyc_C1_div;
  assign T488[52] = cyc_C1_div;
  assign T489[52] = T494[52] | 1'b0;
  assign T489[51] = T494[51] | 1'b0;
  assign T489[50] = T494[50] | 1'b0;
  assign T489[49] = T494[49] | 1'b0;
  assign T489[48] = T494[48] | 1'b0;
  assign T489[47] = T494[47] | 1'b0;
  assign T489[46] = T494[46] | 1'b0;
  assign T489[45] = T494[45] | T928[45];
  assign T489[44] = T494[44] | T928[44];
  assign T489[43] = T494[43] | T928[43];
  assign T489[42] = T494[42] | T928[42];
  assign T489[41] = T494[41] | T928[41];
  assign T489[40] = T494[40] | T928[40];
  assign T489[39] = T494[39] | T928[39];
  assign T489[38] = T494[38] | T928[38];
  assign T489[37] = T494[37] | T928[37];
  assign T489[36] = T494[36] | T928[36];
  assign T489[35] = T494[35] | T928[35];
  assign T489[34] = T494[34] | T928[34];
  assign T489[33] = T494[33] | T928[33];
  assign T489[32] = T494[32] | T928[32];
  assign T489[31] = T494[31] | T928[31];
  assign T489[30] = T494[30] | T928[30];
  assign T489[29] = T494[29] | T928[29];
  assign T489[28] = T494[28] | T928[28];
  assign T489[27] = T494[27] | T928[27];
  assign T489[26] = T494[26] | T928[26];
  assign T489[25] = T494[25] | T928[25];
  assign T489[24] = T494[24] | T928[24];
  assign T489[23] = T494[23] | T928[23];
  assign T489[22] = T494[22] | T928[22];
  assign T489[21] = T494[21] | T928[21];
  assign T489[20] = T494[20] | T928[20];
  assign T489[19] = T494[19] | T928[19];
  assign T489[18] = T494[18] | T928[18];
  assign T489[17] = T494[17] | T928[17];
  assign T489[16] = T494[16] | T928[16];
  assign T489[15] = T494[15] | T928[15];
  assign T489[14] = T494[14] | 1'b0;
  assign T489[13] = T494[13] | 1'b0;
  assign T489[12] = T494[12] | 1'b0;
  assign T489[11] = T494[11] | 1'b0;
  assign T489[10] = T494[10] | 1'b0;
  assign T489[9] = T494[9] | 1'b0;
  assign T489[8] = T494[8] | 1'b0;
  assign T489[7] = T494[7] | 1'b0;
  assign T489[6] = T494[6] | 1'b0;
  assign T489[5] = T494[5] | 1'b0;
  assign T489[4] = T494[4] | 1'b0;
  assign T489[3] = T494[3] | 1'b0;
  assign T489[2] = T494[2] | 1'b0;
  assign T489[1] = T494[1] | 1'b0;
  assign T489[0] = T494[0] | 1'b0;
  assign N152 = ~cyc_C4_sqrt;
  assign cyc_C5_sqrt = N481 & sqrtOp_PB;
  assign T494[52] = T499[52] | 1'b0;
  assign T494[51] = T499[51] | 1'b0;
  assign T494[50] = T499[50] | 1'b0;
  assign T494[49] = T499[49] | 1'b0;
  assign T494[48] = T499[48] | 1'b0;
  assign T494[47] = T499[47] | 1'b0;
  assign T494[46] = T499[46] | 1'b0;
  assign T494[45] = T499[45] | T929[45];
  assign T494[44] = T499[44] | T929[44];
  assign T494[43] = T499[43] | T929[43];
  assign T494[42] = T499[42] | T929[42];
  assign T494[41] = T499[41] | T929[41];
  assign T494[40] = T499[40] | T929[40];
  assign T494[39] = T499[39] | T929[39];
  assign T494[38] = T499[38] | T929[38];
  assign T494[37] = T499[37] | T929[37];
  assign T494[36] = T499[36] | T929[36];
  assign T494[35] = T499[35] | T929[35];
  assign T494[34] = T499[34] | T929[34];
  assign T494[33] = T499[33] | T929[33];
  assign T494[32] = T499[32] | T929[32];
  assign T494[31] = T499[31] | T929[31];
  assign T494[30] = T499[30] | T929[30];
  assign T494[29] = T499[29] | T929[29];
  assign T494[28] = T499[28] | T929[28];
  assign T494[27] = T499[27] | T929[27];
  assign T494[26] = T499[26] | T929[26];
  assign T494[25] = T499[25] | T929[25];
  assign T494[24] = T499[24] | T929[24];
  assign T494[23] = T499[23] | T929[23];
  assign T494[22] = T499[22] | T929[22];
  assign T494[21] = T499[21] | T929[21];
  assign T494[20] = T499[20] | T929[20];
  assign T494[19] = T499[19] | T929[19];
  assign T494[18] = T499[18] | T929[18];
  assign T494[17] = T499[17] | T929[17];
  assign T494[16] = T499[16] | T929[16];
  assign T494[15] = T499[15] | T929[15];
  assign T494[14] = T499[14] | T929[14];
  assign T494[13] = T499[13] | T929[13];
  assign T494[12] = T499[12] | 1'b0;
  assign T494[11] = T499[11] | 1'b0;
  assign T494[10] = T499[10] | 1'b0;
  assign T494[9] = T499[9] | 1'b0;
  assign T494[8] = T499[8] | 1'b0;
  assign T494[7] = T499[7] | 1'b0;
  assign T494[6] = T499[6] | 1'b0;
  assign T494[5] = T499[5] | 1'b0;
  assign T494[4] = T499[4] | 1'b0;
  assign T494[3] = T499[3] | 1'b0;
  assign T494[2] = T499[2] | 1'b0;
  assign T494[1] = T499[1] | 1'b0;
  assign T494[0] = T499[0] | 1'b0;
  assign N153 = ~cyc_C4_div;
  assign cyc_C4_div = N476 & T498;
  assign T498 = ~sqrtOp_PB;
  assign T499[52] = T503[52] | 1'b0;
  assign T499[51] = T503[51] | 1'b0;
  assign T499[50] = T503[50] | 1'b0;
  assign T499[49] = T503[49] | 1'b0;
  assign T499[48] = T503[48] | 1'b0;
  assign T499[47] = T503[47] | 1'b0;
  assign T499[46] = T503[46] | 1'b0;
  assign T499[45] = T503[45] | T930[45];
  assign T499[44] = T503[44] | T930[44];
  assign T499[43] = T503[43] | T930[43];
  assign T499[42] = T503[42] | T930[42];
  assign T499[41] = T503[41] | T930[41];
  assign T499[40] = T503[40] | T930[40];
  assign T499[39] = T503[39] | T930[39];
  assign T499[38] = T503[38] | T930[38];
  assign T499[37] = T503[37] | T930[37];
  assign T499[36] = T503[36] | T930[36];
  assign T499[35] = T503[35] | T930[35];
  assign T499[34] = T503[34] | T930[34];
  assign T499[33] = T503[33] | T930[33];
  assign T499[32] = T503[32] | T930[32];
  assign T499[31] = T503[31] | T930[31];
  assign T499[30] = T503[30] | T930[30];
  assign T499[29] = T503[29] | T930[29];
  assign T499[28] = T503[28] | T930[28];
  assign T499[27] = T503[27] | T930[27];
  assign T499[26] = T503[26] | T930[26];
  assign T499[25] = T503[25] | T930[25];
  assign T499[24] = T503[24] | T930[24];
  assign T499[23] = T503[23] | T930[23];
  assign T499[22] = T503[22] | T930[22];
  assign T499[21] = T503[21] | T930[21];
  assign T499[20] = T503[20] | T930[20];
  assign T499[19] = T503[19] | T930[19];
  assign T499[18] = T503[18] | T930[18];
  assign T499[17] = T503[17] | T930[17];
  assign T499[16] = T503[16] | T930[16];
  assign T499[15] = T503[15] | T930[15];
  assign T499[14] = T503[14] | T930[14];
  assign T499[13] = T503[13] | T930[13];
  assign T499[12] = T503[12] | T930[12];
  assign T499[11] = T503[11] | T930[11];
  assign T499[10] = T503[10] | T930[10];
  assign T499[9] = T503[9] | T930[9];
  assign T499[8] = T503[8] | T930[8];
  assign T499[7] = T503[7] | T930[7];
  assign T499[6] = T503[6] | T930[6];
  assign T499[5] = T503[5] | T930[5];
  assign T499[4] = T503[4] | T930[4];
  assign T499[3] = T503[3] | T930[3];
  assign T499[2] = T503[2] | T930[2];
  assign T499[1] = T503[1] | T930[1];
  assign T499[0] = T503[0] | T930[0];
  assign N154 = ~T502;
  assign T502 = N493 | N308;
  assign T503[52] = T505[52] | 1'b0;
  assign T503[51] = T505[51] | 1'b0;
  assign T503[50] = T505[50] | 1'b0;
  assign T503[49] = T505[49] | 1'b0;
  assign T503[48] = T505[48] | 1'b0;
  assign T503[47] = T505[47] | 1'b0;
  assign T503[46] = T505[46] | 1'b0;
  assign T503[45] = T505[45] | 1'b0;
  assign T503[44] = T505[44] | 1'b0;
  assign T503[43] = T505[43] | 1'b0;
  assign T503[42] = T505[42] | 1'b0;
  assign T503[41] = T505[41] | 1'b0;
  assign T503[40] = T505[40] | 1'b0;
  assign T503[39] = T505[39] | 1'b0;
  assign T503[38] = T505[38] | 1'b0;
  assign T503[37] = T505[37] | 1'b0;
  assign T503[36] = T505[36] | 1'b0;
  assign T503[35] = T505[35] | 1'b0;
  assign T503[34] = T505[34] | 1'b0;
  assign T503[33] = T505[33] | T902[45];
  assign T503[32] = T505[32] | T902[44];
  assign T503[31] = T505[31] | T902[43];
  assign T503[30] = T505[30] | T902[42];
  assign T503[29] = T505[29] | T902[41];
  assign T503[28] = T505[28] | T902[40];
  assign T503[27] = T505[27] | T902[39];
  assign T503[26] = T505[26] | T902[38];
  assign T503[25] = T505[25] | T902[37];
  assign T503[24] = T505[24] | T902[36];
  assign T503[23] = T505[23] | T902[35];
  assign T503[22] = T505[22] | T902[34];
  assign T503[21] = T505[21] | T902[33];
  assign T503[20] = T505[20] | T902[32];
  assign T503[19] = T505[19] | T902[31];
  assign T503[18] = T505[18] | T902[30];
  assign T503[17] = T505[17] | T902[29];
  assign T503[16] = T505[16] | T902[28];
  assign T503[15] = T505[15] | T902[27];
  assign T503[14] = T505[14] | T902[26];
  assign T503[13] = T505[13] | T902[25];
  assign T503[12] = T505[12] | T902[24];
  assign T503[11] = T505[11] | T902[23];
  assign T503[10] = T505[10] | T902[22];
  assign T503[9] = T505[9] | T902[21];
  assign T503[8] = T505[8] | T902[20];
  assign T503[7] = T505[7] | T902[19];
  assign T503[6] = T505[6] | T902[18];
  assign T503[5] = T505[5] | T902[17];
  assign T503[4] = T505[4] | T902[16];
  assign T503[3] = T505[3] | T902[15];
  assign T503[2] = T505[2] | T902[14];
  assign T503[1] = T505[1] | T902[13];
  assign T503[0] = T505[0] | T902[12];
  assign T505[52] = T513[52] | T506[52];
  assign T505[51] = T513[51] | T506[51];
  assign T505[50] = T513[50] | T506[50];
  assign T505[49] = T513[49] | T506[49];
  assign T505[48] = T513[48] | T506[48];
  assign T505[47] = T513[47] | T506[47];
  assign T505[46] = T513[46] | T506[46];
  assign T505[45] = T513[45] | T506[45];
  assign T505[44] = T513[44] | T506[44];
  assign T505[43] = T513[43] | T506[43];
  assign T505[42] = T513[42] | T506[42];
  assign T505[41] = T513[41] | T506[41];
  assign T505[40] = T513[40] | T506[40];
  assign T505[39] = T513[39] | T506[39];
  assign T505[38] = T513[38] | T506[38];
  assign T505[37] = T513[37] | T506[37];
  assign T505[36] = T513[36] | T506[36];
  assign T505[35] = T513[35] | T506[35];
  assign T505[34] = T513[34] | T506[34];
  assign T505[33] = T513[33] | T506[33];
  assign T505[32] = T513[32] | T506[32];
  assign T505[31] = T513[31] | T506[31];
  assign T505[30] = T513[30] | T506[30];
  assign T505[29] = T513[29] | T506[29];
  assign T505[28] = T513[28] | T506[28];
  assign T505[27] = T513[27] | T506[27];
  assign T505[26] = T513[26] | T506[26];
  assign T505[25] = T513[25] | T506[25];
  assign T505[24] = T513[24] | T506[24];
  assign T505[23] = T513[23] | T506[23];
  assign T505[22] = T513[22] | T506[22];
  assign T505[21] = T513[21] | T506[21];
  assign T505[20] = T513[20] | T506[20];
  assign T505[19] = T513[19] | T506[19];
  assign T505[18] = T513[18] | T506[18];
  assign T505[17] = T513[17] | T506[17];
  assign T505[16] = T513[16] | T506[16];
  assign T505[15] = T513[15] | T506[15];
  assign T505[14] = T513[14] | T506[14];
  assign T505[13] = T513[13] | T506[13];
  assign T505[12] = T513[12] | T506[12];
  assign T505[11] = T513[11] | T506[11];
  assign T505[10] = T513[10] | T506[10];
  assign T505[9] = T513[9] | T506[9];
  assign T505[8] = T513[8] | T506[8];
  assign T505[7] = T513[7] | T506[7];
  assign T505[6] = T513[6] | T506[6];
  assign T505[5] = T513[5] | T506[5];
  assign T505[4] = T513[4] | T506[4];
  assign T505[3] = T513[3] | T506[3];
  assign T505[2] = T513[2] | T506[2];
  assign T505[1] = T513[1] | T506[1];
  assign T505[0] = T513[0] | T506[0];
  assign N155 = ~cyc_B6_div;
  assign T506[52] = cyc_B6_div;
  assign cyc_B6_div = T512 & T511;
  assign T511 = ~sqrtOp_PA;
  assign T512 = N502 & valid_PA;
  assign T513[52] = T516[52] | T514[52];
  assign T513[51] = T516[51] | T514[51];
  assign T513[50] = T516[50] | T514[50];
  assign T513[49] = T516[49] | T514[49];
  assign T513[48] = T516[48] | T514[48];
  assign T513[47] = T516[47] | T514[47];
  assign T513[46] = T516[46] | T514[46];
  assign T513[45] = T516[45] | T514[45];
  assign T513[44] = T516[44] | T514[44];
  assign T513[43] = T516[43] | T514[43];
  assign T513[42] = T516[42] | T514[42];
  assign T513[41] = T516[41] | T514[41];
  assign T513[40] = T516[40] | T514[40];
  assign T513[39] = T516[39] | T514[39];
  assign T513[38] = T516[38] | T514[38];
  assign T513[37] = T516[37] | T514[37];
  assign T513[36] = T516[36] | T514[36];
  assign T513[35] = 1'b0 | T514[35];
  assign T513[34] = 1'b0 | T514[34];
  assign T513[33] = 1'b0 | T514[33];
  assign T513[32] = 1'b0 | T514[32];
  assign T513[31] = 1'b0 | T514[31];
  assign T513[30] = 1'b0 | T514[30];
  assign T513[29] = 1'b0 | T514[29];
  assign T513[28] = 1'b0 | T514[28];
  assign T513[27] = 1'b0 | T514[27];
  assign T513[26] = 1'b0 | T514[26];
  assign T513[25] = 1'b0 | T514[25];
  assign T513[24] = 1'b0 | T514[24];
  assign T513[23] = 1'b0 | T514[23];
  assign T513[22] = 1'b0 | T514[22];
  assign T513[21] = 1'b0 | T514[21];
  assign T513[20] = 1'b0 | T514[20];
  assign T513[19] = 1'b0 | T514[19];
  assign T513[18] = 1'b0 | T514[18];
  assign T513[17] = 1'b0 | T514[17];
  assign T513[16] = 1'b0 | T514[16];
  assign T513[15] = 1'b0 | T514[15];
  assign T513[14] = 1'b0 | T514[14];
  assign T513[13] = 1'b0 | T514[13];
  assign T513[12] = 1'b0 | T514[12];
  assign T513[11] = 1'b0 | T514[11];
  assign T513[10] = 1'b0 | T514[10];
  assign T513[9] = 1'b0 | T514[9];
  assign T513[8] = 1'b0 | T514[8];
  assign T513[7] = 1'b0 | T514[7];
  assign T513[6] = 1'b0 | T514[6];
  assign T513[5] = 1'b0 | T514[5];
  assign T513[4] = 1'b0 | T514[4];
  assign T513[3] = 1'b0 | T514[3];
  assign T513[2] = 1'b0 | T514[2];
  assign T513[1] = 1'b0 | T514[1];
  assign T513[0] = 1'b0 | T514[0];
  assign N156 = ~T515;
  assign T514[52] = T515;
  assign T515 = N506 | cyc_A1_div;
  assign io_latchMulAddA_0 = T519 | N312;
  assign T519 = T520 | N476;
  assign T520 = T521 | N308;
  assign T521 = T522 | N493;
  assign T522 = T523 | N513;
  assign T523 = T524 | cyc_B6_div;
  assign T524 = N316 | N506;
  assign io_usingMulAdd[0] = T530 | cyc_B2_sqrt;
  assign cyc_B2_sqrt = N485 & sqrtOp_PB;
  assign T530 = io_latchMulAddA_0 | N502;
  assign io_usingMulAdd[1] = T532 | N285;
  assign T532 = T533 | N481;
  assign T533 = T535 | cyc_B1_sqrt;
  assign cyc_B1_sqrt = N489 & sqrtOp_PB;
  assign T535 = T537 | cyc_B3_sqrt;
  assign cyc_B3_sqrt = N493 & sqrtOp_PB;
  assign T537 = T538 | N513;
  assign T538 = T540 | N498;
  assign T540 = T541 | N506;
  assign T541 = T542 | N294;
  assign T542 = N320 | cyc_A1_div;
  assign io_usingMulAdd[2] = T545 | N509;
  assign T545 = T546 | N308;
  assign T546 = T549 | cyc_B1_div;
  assign cyc_B1_div = N489 & T548;
  assign T548 = ~sqrtOp_PB;
  assign T549 = T550 | cyc_B2_sqrt;
  assign T550 = T553 | cyc_B4_sqrt;
  assign cyc_B4_sqrt = T552 & sqrtOp_PB;
  assign T552 = N513 & valid_PB;
  assign T553 = T554 | N498;
  assign T554 = T555 | N502;
  assign T555 = T556 | N294;
  assign T556 = T558 | N304;
  assign T558 = N330 | cyc_A2_div;
  assign cyc_A2_div = N320 & T559;
  assign T559 = ~sqrtOp_PA;
  assign io_usingMulAdd[3] = T561 | N476;
  assign T561 = T562 | cyc_B1_sqrt;
  assign T562 = T565 | cyc_B2_div;
  assign cyc_B2_div = N485 & T564;
  assign T564 = ~sqrtOp_PB;
  assign T565 = T566 | cyc_B3_sqrt;
  assign T566 = T569 | cyc_B5_sqrt;
  assign cyc_B5_sqrt = T568 & sqrtOp_PB;
  assign T568 = N498 & valid_PB;
  assign T569 = T570 | N502;
  assign T570 = T571 | N506;
  assign T571 = T572 | N304;
  assign T572 = T574 | N299;
  assign T574 = T575 | cyc_A1_div;
  assign T575 = cyc_A4 | cyc_A3_div;
  assign io_exceptionFlags[0] = T705 | T579;
  assign T579 = normalCase_PC & inexactY_E1;
  assign inexactY_E1 = hiRoundPosBit_E1 | anyRoundExtra_E1;
  assign anyRoundExtra_E1 = T676 | T580;
  assign T580 = ~N409;
  assign T581[52] = T673[52] & 1'b0;
  assign T581[51] = T673[51] & T932[51];
  assign T581[50] = T673[50] & T932[50];
  assign T581[49] = T673[49] & T932[49];
  assign T581[48] = T673[48] & T932[48];
  assign T581[47] = T673[47] & T932[47];
  assign T581[46] = T673[46] & T932[46];
  assign T581[45] = T673[45] & T932[45];
  assign T581[44] = T673[44] & T932[44];
  assign T581[43] = T673[43] & T932[43];
  assign T581[42] = T673[42] & T932[42];
  assign T581[41] = T673[41] & T932[41];
  assign T581[40] = T673[40] & T932[40];
  assign T581[39] = T673[39] & T932[39];
  assign T581[38] = T673[38] & T932[38];
  assign T581[37] = T673[37] & T932[37];
  assign T581[36] = T673[36] & T932[36];
  assign T581[35] = T673[35] & T932[35];
  assign T581[34] = T673[34] & T932[34];
  assign T581[33] = T673[33] & T932[33];
  assign T581[32] = T673[32] & T932[32];
  assign T581[31] = T673[31] & T932[31];
  assign T581[30] = T673[30] & T932[30];
  assign T581[29] = T673[29] & T932[29];
  assign T581[28] = T673[28] & T932[28];
  assign T581[27] = T673[27] & T932[27];
  assign T581[26] = T673[26] & T932[26];
  assign T581[25] = T673[25] & T932[25];
  assign T581[24] = T673[24] & T932[24];
  assign T581[23] = T673[23] & T932[23];
  assign T581[22] = T673[22] & T932[22];
  assign T581[21] = T673[21] & T932[21];
  assign T581[20] = T673[20] & T932[20];
  assign T581[19] = T673[19] & T932[19];
  assign T581[18] = T673[18] & T932[18];
  assign T581[17] = T673[17] & T932[17];
  assign T581[16] = T673[16] & T932[16];
  assign T581[15] = T673[15] & T932[15];
  assign T581[14] = T673[14] & T932[14];
  assign T581[13] = T673[13] & T932[13];
  assign T581[12] = T673[12] & T932[12];
  assign T581[11] = T673[11] & T932[11];
  assign T581[10] = T673[10] & T932[10];
  assign T581[9] = T673[9] & T932[9];
  assign T581[8] = T673[8] & T932[8];
  assign T581[7] = T673[7] & T932[7];
  assign T581[6] = T673[6] & T932[6];
  assign T581[5] = T673[5] & T932[5];
  assign T581[4] = T673[4] & T932[4];
  assign T581[3] = T673[3] & T586[0];
  assign T581[2] = T673[2] & T586[1];
  assign T581[1] = T673[1] & T586[2];
  assign T581[0] = T673[0] & T586[3];
  assign T590[12] = ~posExpX_E[12];
  assign T590[11] = ~posExpX_E[11];
  assign T590[10] = ~posExpX_E[10];
  assign T590[9] = ~posExpX_E[9];
  assign T590[8] = ~posExpX_E[8];
  assign T590[7] = ~posExpX_E[7];
  assign T590[6] = ~posExpX_E[6];
  assign T590[5] = ~posExpX_E[5];
  assign T590[4] = ~posExpX_E[4];
  assign T590[3] = ~posExpX_E[3];
  assign T590[2] = ~posExpX_E[2];
  assign T590[1] = ~posExpX_E[1];
  assign T590[0] = ~posExpX_E[0];
  assign sExpX_E[13] = T594[13] | 1'b0;
  assign posExpX_E[12] = T594[12] | T933[12];
  assign posExpX_E[11] = T594[11] | T933[11];
  assign posExpX_E[10] = T594[10] | T933[10];
  assign posExpX_E[9] = T594[9] | T933[9];
  assign posExpX_E[8] = T594[8] | T933[8];
  assign posExpX_E[7] = T594[7] | T933[7];
  assign posExpX_E[6] = T594[6] | T933[6];
  assign posExpX_E[5] = T594[5] | T933[5];
  assign posExpX_E[4] = T594[4] | T933[4];
  assign posExpX_E[3] = T594[3] | T933[3];
  assign posExpX_E[2] = T594[2] | T933[2];
  assign posExpX_E[1] = T594[1] | T933[1];
  assign posExpX_E[0] = T594[0] | T933[0];
  assign T594[13] = T604[13] | T595[13];
  assign T594[12] = T604[12] | T595[12];
  assign T594[11] = T604[11] | T595[11];
  assign T594[10] = T604[10] | T595[10];
  assign T594[9] = T604[9] | T595[9];
  assign T594[8] = T604[8] | T595[8];
  assign T594[7] = T604[7] | T595[7];
  assign T594[6] = T604[6] | T595[6];
  assign T594[5] = T604[5] | T595[5];
  assign T594[4] = T604[4] | T595[4];
  assign T594[3] = T604[3] | T595[3];
  assign T594[2] = T604[2] | T595[2];
  assign T594[1] = T604[1] | T595[1];
  assign T594[0] = T604[0] | T595[0];
  assign N157 = ~T601;
  assign expP1_PC[0] = N130;
  assign T601 = T603 & T602;
  assign T602 = ~E_E_div;
  assign T603 = ~sqrtOp_PC;
  assign N158 = ~T605;
  assign T605 = T606 & E_E_div;
  assign T606 = ~sqrtOp_PC;
  assign T932[19] = 1'b0 | T618[15];
  assign T932[18] = T621[15] | 1'b0;
  assign T932[17] = 1'b0 | T618_13;
  assign T932[16] = T619[14] | 1'b0;
  assign T932[15] = 1'b0 | T618_11;
  assign T932[14] = T619_12 | 1'b0;
  assign T932[13] = 1'b0 | T618_9;
  assign T932[12] = T619_10 | 1'b0;
  assign T932[11] = 1'b0 | T618_7;
  assign T932[10] = T619_8 | 1'b0;
  assign T932[9] = 1'b0 | T618_5;
  assign T932[8] = T619_6 | 1'b0;
  assign T932[7] = 1'b0 | T618_3;
  assign T932[6] = T619_4 | 1'b0;
  assign T932[5] = 1'b0 | T618_1;
  assign T932[4] = T619_2 | 1'b0;
  assign T621[15] = 1'b0 | T622[15];
  assign T618[15] = 1'b0 | T622[14];
  assign T619[14] = T625[15] | 1'b0;
  assign T618_13 = T625[14] | 1'b0;
  assign T619_12 = 1'b0 | T622_11;
  assign T618_11 = 1'b0 | T622_10;
  assign T619_10 = T623[13] | 1'b0;
  assign T618_9 = T623[12] | 1'b0;
  assign T619_8 = 1'b0 | T622_7;
  assign T618_7 = 1'b0 | T622_6;
  assign T619_6 = T623_9 | 1'b0;
  assign T618_5 = T623_8 | 1'b0;
  assign T619_4 = 1'b0 | T622_3;
  assign T618_3 = 1'b0 | T622_2;
  assign T619_2 = T623_5 | 1'b0;
  assign T618_1 = T623_4 | 1'b0;
  assign T625[15] = 1'b0 | T626[15];
  assign T625[14] = 1'b0 | T626[14];
  assign T622[15] = 1'b0 | T626[13];
  assign T622[14] = 1'b0 | T626[12];
  assign T623[13] = T629[15] | 1'b0;
  assign T623[12] = T629[14] | 1'b0;
  assign T622_11 = T629[13] | 1'b0;
  assign T622_10 = T629[12] | 1'b0;
  assign T623_9 = 1'b0 | T626_7;
  assign T623_8 = 1'b0 | T626_6;
  assign T622_7 = 1'b0 | T626_5;
  assign T622_6 = 1'b0 | T626_4;
  assign T623_5 = T627[11] | 1'b0;
  assign T623_4 = T627[10] | 1'b0;
  assign T622_3 = T627[9] | 1'b0;
  assign T622_2 = T627[8] | 1'b0;
  assign T629[15] = 1'b0 | T587[7];
  assign T629[14] = 1'b0 | T587[6];
  assign T629[13] = 1'b0 | T587[5];
  assign T629[12] = 1'b0 | T587[4];
  assign T626[15] = 1'b0 | T587[3];
  assign T626[14] = 1'b0 | T587[2];
  assign T626[13] = 1'b0 | T587[1];
  assign T626[12] = 1'b0 | T587[0];
  assign T627[11] = T587[15] | 1'b0;
  assign T627[10] = T587[14] | 1'b0;
  assign T627[9] = T587[13] | 1'b0;
  assign T627[8] = T587[12] | 1'b0;
  assign T626_7 = T587[11] | 1'b0;
  assign T626_6 = T587[10] | 1'b0;
  assign T626_5 = T587[9] | 1'b0;
  assign T626_4 = T587[8] | 1'b0;
  assign T932[51] = 1'b0 | T643[31];
  assign T932[50] = T646[31] | 1'b0;
  assign T932[49] = 1'b0 | T643_29;
  assign T932[48] = T644[30] | 1'b0;
  assign T932[47] = 1'b0 | T643_27;
  assign T932[46] = T644_28 | 1'b0;
  assign T932[45] = 1'b0 | T643_25;
  assign T932[44] = T644_26 | 1'b0;
  assign T932[43] = 1'b0 | T643_23;
  assign T932[42] = T644_24 | 1'b0;
  assign T932[41] = 1'b0 | T643_21;
  assign T932[40] = T644_22 | 1'b0;
  assign T932[39] = 1'b0 | T643_19;
  assign T932[38] = T644_20 | 1'b0;
  assign T932[37] = 1'b0 | T643_17;
  assign T932[36] = T644_18 | 1'b0;
  assign T932[35] = 1'b0 | T643_15;
  assign T932[34] = T644_16 | 1'b0;
  assign T932[33] = 1'b0 | T643_13;
  assign T932[32] = T644_14 | 1'b0;
  assign T932[31] = 1'b0 | T643_11;
  assign T932[30] = T644_12 | 1'b0;
  assign T932[29] = 1'b0 | T643_9;
  assign T932[28] = T644_10 | 1'b0;
  assign T932[27] = 1'b0 | T643_7;
  assign T932[26] = T644_8 | 1'b0;
  assign T932[25] = 1'b0 | T643_5;
  assign T932[24] = T644_6 | 1'b0;
  assign T932[23] = 1'b0 | T643_3;
  assign T932[22] = T644_4 | 1'b0;
  assign T932[21] = 1'b0 | T643_1;
  assign T932[20] = T644_2 | 1'b0;
  assign T646[31] = 1'b0 | T647[31];
  assign T643[31] = 1'b0 | T647[30];
  assign T644[30] = T650[31] | 1'b0;
  assign T643_29 = T650[30] | 1'b0;
  assign T644_28 = 1'b0 | T647_27;
  assign T643_27 = 1'b0 | T647_26;
  assign T644_26 = T648[29] | 1'b0;
  assign T643_25 = T648[28] | 1'b0;
  assign T644_24 = 1'b0 | T647_23;
  assign T643_23 = 1'b0 | T647_22;
  assign T644_22 = T648_25 | 1'b0;
  assign T643_21 = T648_24 | 1'b0;
  assign T644_20 = 1'b0 | T647_19;
  assign T643_19 = 1'b0 | T647_18;
  assign T644_18 = T648_21 | 1'b0;
  assign T643_17 = T648_20 | 1'b0;
  assign T644_16 = 1'b0 | T647_15;
  assign T643_15 = 1'b0 | T647_14;
  assign T644_14 = T648_17 | 1'b0;
  assign T643_13 = T648_16 | 1'b0;
  assign T644_12 = 1'b0 | T647_11;
  assign T643_11 = 1'b0 | T647_10;
  assign T644_10 = T648_13 | 1'b0;
  assign T643_9 = T648_12 | 1'b0;
  assign T644_8 = 1'b0 | T647_7;
  assign T643_7 = 1'b0 | T647_6;
  assign T644_6 = T648_9 | 1'b0;
  assign T643_5 = T648_8 | 1'b0;
  assign T644_4 = 1'b0 | T647_3;
  assign T643_3 = 1'b0 | T647_2;
  assign T644_2 = T648_5 | 1'b0;
  assign T643_1 = T648_4 | 1'b0;
  assign T650[31] = 1'b0 | T651[31];
  assign T650[30] = 1'b0 | T651[30];
  assign T647[31] = 1'b0 | T651[29];
  assign T647[30] = 1'b0 | T651[28];
  assign T648[29] = T654[31] | 1'b0;
  assign T648[28] = T654[30] | 1'b0;
  assign T647_27 = T654[29] | 1'b0;
  assign T647_26 = T654[28] | 1'b0;
  assign T648_25 = 1'b0 | T651_23;
  assign T648_24 = 1'b0 | T651_22;
  assign T647_23 = 1'b0 | T651_21;
  assign T647_22 = 1'b0 | T651_20;
  assign T648_21 = T652[27] | 1'b0;
  assign T648_20 = T652[26] | 1'b0;
  assign T647_19 = T652[25] | 1'b0;
  assign T647_18 = T652[24] | 1'b0;
  assign T648_17 = 1'b0 | T651_15;
  assign T648_16 = 1'b0 | T651_14;
  assign T647_15 = 1'b0 | T651_13;
  assign T647_14 = 1'b0 | T651_12;
  assign T648_13 = T652_19 | 1'b0;
  assign T648_12 = T652_18 | 1'b0;
  assign T647_11 = T652_17 | 1'b0;
  assign T647_10 = T652_16 | 1'b0;
  assign T648_9 = 1'b0 | T651_7;
  assign T648_8 = 1'b0 | T651_6;
  assign T647_7 = 1'b0 | T651_5;
  assign T647_6 = 1'b0 | T651_4;
  assign T648_5 = T652_11 | 1'b0;
  assign T648_4 = T652_10 | 1'b0;
  assign T647_3 = T652_9 | 1'b0;
  assign T647_2 = T652_8 | 1'b0;
  assign T654[31] = 1'b0 | T655[31];
  assign T654[30] = 1'b0 | T655[30];
  assign T654[29] = 1'b0 | T655[29];
  assign T654[28] = 1'b0 | T655[28];
  assign T651[31] = 1'b0 | T655[27];
  assign T651[30] = 1'b0 | T655[26];
  assign T651[29] = 1'b0 | T655[25];
  assign T651[28] = 1'b0 | T655[24];
  assign T652[27] = T658[31] | 1'b0;
  assign T652[26] = T658[30] | 1'b0;
  assign T652[25] = T658[29] | 1'b0;
  assign T652[24] = T658[28] | 1'b0;
  assign T651_23 = T658[27] | 1'b0;
  assign T651_22 = T658[26] | 1'b0;
  assign T651_21 = T658[25] | 1'b0;
  assign T651_20 = T658[24] | 1'b0;
  assign T652_19 = 1'b0 | T655_15;
  assign T652_18 = 1'b0 | T655_14;
  assign T652_17 = 1'b0 | T655_13;
  assign T652_16 = 1'b0 | T655_12;
  assign T651_15 = 1'b0 | T655_11;
  assign T651_14 = 1'b0 | T655_10;
  assign T651_13 = 1'b0 | T655_9;
  assign T651_12 = 1'b0 | T655_8;
  assign T652_11 = T656[23] | 1'b0;
  assign T652_10 = T656[22] | 1'b0;
  assign T652_9 = T656[21] | 1'b0;
  assign T652_8 = T656[20] | 1'b0;
  assign T651_7 = T656[19] | 1'b0;
  assign T651_6 = T656[18] | 1'b0;
  assign T651_5 = T656[17] | 1'b0;
  assign T651_4 = T656[16] | 1'b0;
  assign T658[31] = 1'b0 | T588[15];
  assign T658[30] = 1'b0 | T588[14];
  assign T658[29] = 1'b0 | T588[13];
  assign T658[28] = 1'b0 | T588[12];
  assign T658[27] = 1'b0 | T588[11];
  assign T658[26] = 1'b0 | T588[10];
  assign T658[25] = 1'b0 | T588[9];
  assign T658[24] = 1'b0 | T588[8];
  assign T655[31] = 1'b0 | T588[7];
  assign T655[30] = 1'b0 | T588[6];
  assign T655[29] = 1'b0 | T588[5];
  assign T655[28] = 1'b0 | T588[4];
  assign T655[27] = 1'b0 | T588[3];
  assign T655[26] = 1'b0 | T588[2];
  assign T655[25] = 1'b0 | T588[1];
  assign T655[24] = 1'b0 | T588[0];
  assign T656[23] = T588[31] | 1'b0;
  assign T656[22] = T588[30] | 1'b0;
  assign T656[21] = T588[29] | 1'b0;
  assign T656[20] = T588[28] | 1'b0;
  assign T656[19] = T588[27] | 1'b0;
  assign T656[18] = T588[26] | 1'b0;
  assign T656[17] = T588[25] | 1'b0;
  assign T656[16] = T588[24] | 1'b0;
  assign T655_15 = T588[23] | 1'b0;
  assign T655_14 = T588[22] | 1'b0;
  assign T655_13 = T588[21] | 1'b0;
  assign T655_12 = T588[20] | 1'b0;
  assign T655_11 = T588[19] | 1'b0;
  assign T655_10 = T588[18] | 1'b0;
  assign T655_9 = T588[17] | 1'b0;
  assign T655_8 = T588[16] | 1'b0;
  assign T673[52] = ~T727[52];
  assign T673[51] = ~T727[51];
  assign T673[50] = ~T727[50];
  assign T673[49] = ~T727[49];
  assign T673[48] = ~T727[48];
  assign T673[47] = ~T727[47];
  assign T673[46] = ~T727[46];
  assign T673[45] = ~T727[45];
  assign T673[44] = ~T727[44];
  assign T673[43] = ~T727[43];
  assign T673[42] = ~T727[42];
  assign T673[41] = ~T727[41];
  assign T673[40] = ~T727[40];
  assign T673[39] = ~T727[39];
  assign T673[38] = ~T727[38];
  assign T673[37] = ~T727[37];
  assign T673[36] = ~T727[36];
  assign T673[35] = ~T727[35];
  assign T673[34] = ~T727[34];
  assign T673[33] = ~T727[33];
  assign T673[32] = ~T727[32];
  assign T673[31] = ~T727[31];
  assign T673[30] = ~T727[30];
  assign T673[29] = ~T727[29];
  assign T673[28] = ~T727[28];
  assign T673[27] = ~T727[27];
  assign T673[26] = ~T727[26];
  assign T673[25] = ~T727[25];
  assign T673[24] = ~T727[24];
  assign T673[23] = ~T727[23];
  assign T673[22] = ~T727[22];
  assign T673[21] = ~T727[21];
  assign T673[20] = ~T727[20];
  assign T673[19] = ~T727[19];
  assign T673[18] = ~T727[18];
  assign T673[17] = ~T727[17];
  assign T673[16] = ~T727[16];
  assign T673[15] = ~T727[15];
  assign T673[14] = ~T727[14];
  assign T673[13] = ~T727[13];
  assign T673[12] = ~T727[12];
  assign T673[11] = ~T727[11];
  assign T673[10] = ~T727[10];
  assign T673[9] = ~T727[9];
  assign T673[8] = ~T727[8];
  assign T673[7] = ~T727[7];
  assign T673[6] = ~T727[6];
  assign T673[5] = ~T727[5];
  assign T673[4] = ~T727[4];
  assign T673[3] = ~T727[3];
  assign T673[2] = ~T727[2];
  assign T673[1] = ~T727[1];
  assign T673[0] = ~T727[0];
  assign T676 = T678 | T677;
  assign T677 = ~extraT_E;
  assign T678 = ~isZeroRemT_E;
  assign T680 = N266 & T681;
  assign T681 = T684 | N268;
  assign T684 = ~sqrtOp_PC;
  assign hiRoundPosBit_E1 = N463 ^ T688;
  assign T688 = T689 & extraT_E;
  assign T689 = T690 & N409;
  assign T690 = roundMask_E[0] & T691;
  assign T691 = ~trueLtX_E1;
  assign T696 = T698 & T697;
  assign T697 = ~isZeroRemT_E;
  assign T698 = ~isNegRemT_E;
  assign T700[52] = T727[52] & T701[52];
  assign T700[51] = T727[51] & T701[51];
  assign T700[50] = T727[50] & T701[50];
  assign T700[49] = T727[49] & T701[49];
  assign T700[48] = T727[48] & T701[48];
  assign T700[47] = T727[47] & T701[47];
  assign T700[46] = T727[46] & T701[46];
  assign T700[45] = T727[45] & T701[45];
  assign T700[44] = T727[44] & T701[44];
  assign T700[43] = T727[43] & T701[43];
  assign T700[42] = T727[42] & T701[42];
  assign T700[41] = T727[41] & T701[41];
  assign T700[40] = T727[40] & T701[40];
  assign T700[39] = T727[39] & T701[39];
  assign T700[38] = T727[38] & T701[38];
  assign T700[37] = T727[37] & T701[37];
  assign T700[36] = T727[36] & T701[36];
  assign T700[35] = T727[35] & T701[35];
  assign T700[34] = T727[34] & T701[34];
  assign T700[33] = T727[33] & T701[33];
  assign T700[32] = T727[32] & T701[32];
  assign T700[31] = T727[31] & T701[31];
  assign T700[30] = T727[30] & T701[30];
  assign T700[29] = T727[29] & T701[29];
  assign T700[28] = T727[28] & T701[28];
  assign T700[27] = T727[27] & T701[27];
  assign T700[26] = T727[26] & T701[26];
  assign T700[25] = T727[25] & T701[25];
  assign T700[24] = T727[24] & T701[24];
  assign T700[23] = T727[23] & T701[23];
  assign T700[22] = T727[22] & T701[22];
  assign T700[21] = T727[21] & T701[21];
  assign T700[20] = T727[20] & T701[20];
  assign T700[19] = T727[19] & T701[19];
  assign T700[18] = T727[18] & T701[18];
  assign T700[17] = T727[17] & T701[17];
  assign T700[16] = T727[16] & T701[16];
  assign T700[15] = T727[15] & T701[15];
  assign T700[14] = T727[14] & T701[14];
  assign T700[13] = T727[13] & T701[13];
  assign T700[12] = T727[12] & T701[12];
  assign T700[11] = T727[11] & T701[11];
  assign T700[10] = T727[10] & T701[10];
  assign T700[9] = T727[9] & T701[9];
  assign T700[8] = T727[8] & T701[8];
  assign T700[7] = T727[7] & T701[7];
  assign T700[6] = T727[6] & T701[6];
  assign T700[5] = T727[5] & T701[5];
  assign T700[4] = T727[4] & T701[4];
  assign T700[3] = T727[3] & T701[3];
  assign T700[2] = T727[2] & T701[2];
  assign T700[1] = T727[1] & T701[1];
  assign T700[0] = T727[0] & T701[0];
  assign T701[52] = T703[53] & T932[51];
  assign T701[51] = T703[52] & T932[50];
  assign T701[50] = T703[51] & T932[49];
  assign T701[49] = T703[50] & T932[48];
  assign T701[48] = T703[49] & T932[47];
  assign T701[47] = T703[48] & T932[46];
  assign T701[46] = T703[47] & T932[45];
  assign T701[45] = T703[46] & T932[44];
  assign T701[44] = T703[45] & T932[43];
  assign T701[43] = T703[44] & T932[42];
  assign T701[42] = T703[43] & T932[41];
  assign T701[41] = T703[42] & T932[40];
  assign T701[40] = T703[41] & T932[39];
  assign T701[39] = T703[40] & T932[38];
  assign T701[38] = T703[39] & T932[37];
  assign T701[37] = T703[38] & T932[36];
  assign T701[36] = T703[37] & T932[35];
  assign T701[35] = T703[36] & T932[34];
  assign T701[34] = T703[35] & T932[33];
  assign T701[33] = T703[34] & T932[32];
  assign T701[32] = T703[33] & T932[31];
  assign T701[31] = T703[32] & T932[30];
  assign T701[30] = T703[31] & T932[29];
  assign T701[29] = T703[30] & T932[28];
  assign T701[28] = T703[29] & T932[27];
  assign T701[27] = T703[28] & T932[26];
  assign T701[26] = T703[27] & T932[25];
  assign T701[25] = T703[26] & T932[24];
  assign T701[24] = T703[25] & T932[23];
  assign T701[23] = T703[24] & T932[22];
  assign T701[22] = T703[23] & T932[21];
  assign T701[21] = T703[22] & T932[20];
  assign T701[20] = T703[21] & T932[19];
  assign T701[19] = T703[20] & T932[18];
  assign T701[18] = T703[19] & T932[17];
  assign T701[17] = T703[18] & T932[16];
  assign T701[16] = T703[17] & T932[15];
  assign T701[15] = T703[16] & T932[14];
  assign T701[14] = T703[15] & T932[13];
  assign T701[13] = T703[14] & T932[12];
  assign T701[12] = T703[13] & T932[11];
  assign T701[11] = T703[12] & T932[10];
  assign T701[10] = T703[11] & T932[9];
  assign T701[9] = T703[10] & T932[8];
  assign T701[8] = T703[9] & T932[7];
  assign T701[7] = T703[8] & T932[6];
  assign T701[6] = T703[7] & T932[5];
  assign T701[5] = T703[6] & T932[4];
  assign T701[4] = T703[5] & T586[0];
  assign T701[3] = T703[4] & T586[1];
  assign T701[2] = T703[3] & T586[2];
  assign T701[1] = T703[2] & T586[3];
  assign T701[0] = T703[1] & roundMask_E[0];
  assign incrPosMask_E[0] = T703[0] & 1'b1;
  assign T703[53] = ~1'b0;
  assign T703[52] = ~T932[51];
  assign T703[51] = ~T932[50];
  assign T703[50] = ~T932[49];
  assign T703[49] = ~T932[48];
  assign T703[48] = ~T932[47];
  assign T703[47] = ~T932[46];
  assign T703[46] = ~T932[45];
  assign T703[45] = ~T932[44];
  assign T703[44] = ~T932[43];
  assign T703[43] = ~T932[42];
  assign T703[42] = ~T932[41];
  assign T703[41] = ~T932[40];
  assign T703[40] = ~T932[39];
  assign T703[39] = ~T932[38];
  assign T703[38] = ~T932[37];
  assign T703[37] = ~T932[36];
  assign T703[36] = ~T932[35];
  assign T703[35] = ~T932[34];
  assign T703[34] = ~T932[33];
  assign T703[33] = ~T932[32];
  assign T703[32] = ~T932[31];
  assign T703[31] = ~T932[30];
  assign T703[30] = ~T932[29];
  assign T703[29] = ~T932[28];
  assign T703[28] = ~T932[27];
  assign T703[27] = ~T932[26];
  assign T703[26] = ~T932[25];
  assign T703[25] = ~T932[24];
  assign T703[24] = ~T932[23];
  assign T703[23] = ~T932[22];
  assign T703[22] = ~T932[21];
  assign T703[21] = ~T932[20];
  assign T703[20] = ~T932[19];
  assign T703[19] = ~T932[18];
  assign T703[18] = ~T932[17];
  assign T703[17] = ~T932[16];
  assign T703[16] = ~T932[15];
  assign T703[15] = ~T932[14];
  assign T703[14] = ~T932[13];
  assign T703[13] = ~T932[12];
  assign T703[12] = ~T932[11];
  assign T703[11] = ~T932[10];
  assign T703[10] = ~T932[9];
  assign T703[9] = ~T932[8];
  assign T703[8] = ~T932[7];
  assign T703[7] = ~T932[6];
  assign T703[6] = ~T932[5];
  assign T703[5] = ~T932[4];
  assign T703[4] = ~T586[0];
  assign T703[3] = ~T586[1];
  assign T703[2] = ~T586[2];
  assign T703[1] = ~T586[3];
  assign T703[0] = ~roundMask_E[0];
  assign T705 = io_exceptionFlags[2] | io_exceptionFlags[1];
  assign io_exceptionFlags[1] = normalCase_PC & underflowY_E1;
  assign underflowY_E1 = totalUnderflowY_E1 | T706;
  assign T706 = T707 & inexactY_E1;
  assign totalUnderflowY_E1 = sExpY_E1[13] | T708;
  assign sExpY_E1[13] = T759[13] | 1'b0;
  assign T709[12] = T759[12] | T943[12];
  assign T709[11] = T759[11] | T943[11];
  assign T709[10] = T759[10] | T943[10];
  assign T709[9] = T759[9] | T943[9];
  assign T709[8] = T759[8] | T943[8];
  assign T709[7] = T759[7] | T943[7];
  assign T709[6] = T759[6] | T943[6];
  assign T709[5] = T759[5] | T943[5];
  assign T709[4] = T759[4] | T943[4];
  assign T709[3] = T759[3] | T943[3];
  assign T709[2] = T759[2] | T943[2];
  assign T709[1] = T759[1] | T943[1];
  assign T709[0] = T759[0] | T943[0];
  assign N159 = ~T713;
  assign T713 = sigY_E1_53 & sqrtOp_PC;
  assign sigY_E1_53 = T724_53 & T715_53;
  assign sigY_E1[51] = T724[51] & T715[51];
  assign sigY_E1[50] = T724[50] & T715[50];
  assign sigY_E1[49] = T724[49] & T715[49];
  assign sigY_E1[48] = T724[48] & T715[48];
  assign sigY_E1[47] = T724[47] & T715[47];
  assign sigY_E1[46] = T724[46] & T715[46];
  assign sigY_E1[45] = T724[45] & T715[45];
  assign sigY_E1[44] = T724[44] & T715[44];
  assign sigY_E1[43] = T724[43] & T715[43];
  assign sigY_E1[42] = T724[42] & T715[42];
  assign sigY_E1[41] = T724[41] & T715[41];
  assign sigY_E1[40] = T724[40] & T715[40];
  assign sigY_E1[39] = T724[39] & T715[39];
  assign sigY_E1[38] = T724[38] & T715[38];
  assign sigY_E1[37] = T724[37] & T715[37];
  assign sigY_E1[36] = T724[36] & T715[36];
  assign sigY_E1[35] = T724[35] & T715[35];
  assign sigY_E1[34] = T724[34] & T715[34];
  assign sigY_E1[33] = T724[33] & T715[33];
  assign sigY_E1[32] = T724[32] & T715[32];
  assign sigY_E1[31] = T724[31] & T715[31];
  assign sigY_E1[30] = T724[30] & T715[30];
  assign sigY_E1[29] = T724[29] & T715[29];
  assign sigY_E1[28] = T724[28] & T715[28];
  assign sigY_E1[27] = T724[27] & T715[27];
  assign sigY_E1[26] = T724[26] & T715[26];
  assign sigY_E1[25] = T724[25] & T715[25];
  assign sigY_E1[24] = T724[24] & T715[24];
  assign sigY_E1[23] = T724[23] & T715[23];
  assign sigY_E1[22] = T724[22] & T715[22];
  assign sigY_E1[21] = T724[21] & T715[21];
  assign sigY_E1[20] = T724[20] & T715[20];
  assign sigY_E1[19] = T724[19] & T715[19];
  assign sigY_E1[18] = T724[18] & T715[18];
  assign sigY_E1[17] = T724[17] & T715[17];
  assign sigY_E1[16] = T724[16] & T715[16];
  assign sigY_E1[15] = T724[15] & T715[15];
  assign sigY_E1[14] = T724[14] & T715[14];
  assign sigY_E1[13] = T724[13] & T715[13];
  assign sigY_E1[12] = T724[12] & T715[12];
  assign sigY_E1[11] = T724[11] & T715[11];
  assign sigY_E1[10] = T724[10] & T715[10];
  assign sigY_E1[9] = T724[9] & T715[9];
  assign sigY_E1[8] = T724[8] & T715[8];
  assign sigY_E1[7] = T724[7] & T715[7];
  assign sigY_E1[6] = T724[6] & T715[6];
  assign sigY_E1[5] = T724[5] & T715[5];
  assign sigY_E1[4] = T724[4] & T715[4];
  assign sigY_E1[3] = T724[3] & T715[3];
  assign sigY_E1[2] = T724[2] & T715[2];
  assign sigY_E1[1] = T724[1] & T715[1];
  assign sigY_E1[0] = T724[0] & T715[0];
  assign T715_53 = ~roundEvenMask_E1_53;
  assign T715[51] = ~roundEvenMask_E1[51];
  assign T715[50] = ~roundEvenMask_E1[50];
  assign T715[49] = ~roundEvenMask_E1[49];
  assign T715[48] = ~roundEvenMask_E1[48];
  assign T715[47] = ~roundEvenMask_E1[47];
  assign T715[46] = ~roundEvenMask_E1[46];
  assign T715[45] = ~roundEvenMask_E1[45];
  assign T715[44] = ~roundEvenMask_E1[44];
  assign T715[43] = ~roundEvenMask_E1[43];
  assign T715[42] = ~roundEvenMask_E1[42];
  assign T715[41] = ~roundEvenMask_E1[41];
  assign T715[40] = ~roundEvenMask_E1[40];
  assign T715[39] = ~roundEvenMask_E1[39];
  assign T715[38] = ~roundEvenMask_E1[38];
  assign T715[37] = ~roundEvenMask_E1[37];
  assign T715[36] = ~roundEvenMask_E1[36];
  assign T715[35] = ~roundEvenMask_E1[35];
  assign T715[34] = ~roundEvenMask_E1[34];
  assign T715[33] = ~roundEvenMask_E1[33];
  assign T715[32] = ~roundEvenMask_E1[32];
  assign T715[31] = ~roundEvenMask_E1[31];
  assign T715[30] = ~roundEvenMask_E1[30];
  assign T715[29] = ~roundEvenMask_E1[29];
  assign T715[28] = ~roundEvenMask_E1[28];
  assign T715[27] = ~roundEvenMask_E1[27];
  assign T715[26] = ~roundEvenMask_E1[26];
  assign T715[25] = ~roundEvenMask_E1[25];
  assign T715[24] = ~roundEvenMask_E1[24];
  assign T715[23] = ~roundEvenMask_E1[23];
  assign T715[22] = ~roundEvenMask_E1[22];
  assign T715[21] = ~roundEvenMask_E1[21];
  assign T715[20] = ~roundEvenMask_E1[20];
  assign T715[19] = ~roundEvenMask_E1[19];
  assign T715[18] = ~roundEvenMask_E1[18];
  assign T715[17] = ~roundEvenMask_E1[17];
  assign T715[16] = ~roundEvenMask_E1[16];
  assign T715[15] = ~roundEvenMask_E1[15];
  assign T715[14] = ~roundEvenMask_E1[14];
  assign T715[13] = ~roundEvenMask_E1[13];
  assign T715[12] = ~roundEvenMask_E1[12];
  assign T715[11] = ~roundEvenMask_E1[11];
  assign T715[10] = ~roundEvenMask_E1[10];
  assign T715[9] = ~roundEvenMask_E1[9];
  assign T715[8] = ~roundEvenMask_E1[8];
  assign T715[7] = ~roundEvenMask_E1[7];
  assign T715[6] = ~roundEvenMask_E1[6];
  assign T715[5] = ~roundEvenMask_E1[5];
  assign T715[4] = ~roundEvenMask_E1[4];
  assign T715[3] = ~roundEvenMask_E1[3];
  assign T715[2] = ~roundEvenMask_E1[2];
  assign T715[1] = ~roundEvenMask_E1[1];
  assign T715[0] = ~roundEvenMask_E1[0];
  assign N160 = ~T716;
  assign T716 = T718 & T717;
  assign T717 = ~anyRoundExtra_E1;
  assign T718 = N411 & hiRoundPosBit_E1;
  assign N161 = ~T730;
  assign sigY0_E_53 = sigAdjT_E[53] & 1'b1;
  assign sigY0_E[51] = sigAdjT_E[51] & T725[51];
  assign sigY0_E[50] = sigAdjT_E[50] & T725[50];
  assign sigY0_E[49] = sigAdjT_E[49] & T725[49];
  assign sigY0_E[48] = sigAdjT_E[48] & T725[48];
  assign sigY0_E[47] = sigAdjT_E[47] & T725[47];
  assign sigY0_E[46] = sigAdjT_E[46] & T725[46];
  assign sigY0_E[45] = sigAdjT_E[45] & T725[45];
  assign sigY0_E[44] = sigAdjT_E[44] & T725[44];
  assign sigY0_E[43] = sigAdjT_E[43] & T725[43];
  assign sigY0_E[42] = sigAdjT_E[42] & T725[42];
  assign sigY0_E[41] = sigAdjT_E[41] & T725[41];
  assign sigY0_E[40] = sigAdjT_E[40] & T725[40];
  assign sigY0_E[39] = sigAdjT_E[39] & T725[39];
  assign sigY0_E[38] = sigAdjT_E[38] & T725[38];
  assign sigY0_E[37] = sigAdjT_E[37] & T725[37];
  assign sigY0_E[36] = sigAdjT_E[36] & T725[36];
  assign sigY0_E[35] = sigAdjT_E[35] & T725[35];
  assign sigY0_E[34] = sigAdjT_E[34] & T725[34];
  assign sigY0_E[33] = sigAdjT_E[33] & T725[33];
  assign sigY0_E[32] = sigAdjT_E[32] & T725[32];
  assign sigY0_E[31] = sigAdjT_E[31] & T725[31];
  assign sigY0_E[30] = sigAdjT_E[30] & T725[30];
  assign sigY0_E[29] = sigAdjT_E[29] & T725[29];
  assign sigY0_E[28] = sigAdjT_E[28] & T725[28];
  assign sigY0_E[27] = sigAdjT_E[27] & T725[27];
  assign sigY0_E[26] = sigAdjT_E[26] & T725[26];
  assign sigY0_E[25] = sigAdjT_E[25] & T725[25];
  assign sigY0_E[24] = sigAdjT_E[24] & T725[24];
  assign sigY0_E[23] = sigAdjT_E[23] & T725[23];
  assign sigY0_E[22] = sigAdjT_E[22] & T725[22];
  assign sigY0_E[21] = sigAdjT_E[21] & T725[21];
  assign sigY0_E[20] = sigAdjT_E[20] & T725[20];
  assign sigY0_E[19] = sigAdjT_E[19] & T725[19];
  assign sigY0_E[18] = sigAdjT_E[18] & T725[18];
  assign sigY0_E[17] = sigAdjT_E[17] & T725[17];
  assign sigY0_E[16] = sigAdjT_E[16] & T725[16];
  assign sigY0_E[15] = sigAdjT_E[15] & T725[15];
  assign sigY0_E[14] = sigAdjT_E[14] & T725[14];
  assign sigY0_E[13] = sigAdjT_E[13] & T725[13];
  assign sigY0_E[12] = sigAdjT_E[12] & T725[12];
  assign sigY0_E[11] = sigAdjT_E[11] & T725[11];
  assign sigY0_E[10] = sigAdjT_E[10] & T725[10];
  assign sigY0_E[9] = sigAdjT_E[9] & T725[9];
  assign sigY0_E[8] = sigAdjT_E[8] & T725[8];
  assign sigY0_E[7] = sigAdjT_E[7] & T725[7];
  assign sigY0_E[6] = sigAdjT_E[6] & T725[6];
  assign sigY0_E[5] = sigAdjT_E[5] & T725[5];
  assign sigY0_E[4] = sigAdjT_E[4] & T725[4];
  assign sigY0_E[3] = sigAdjT_E[3] & T725[3];
  assign sigY0_E[2] = sigAdjT_E[2] & T725[2];
  assign sigY0_E[1] = sigAdjT_E[1] & T725[1];
  assign sigY0_E[0] = sigAdjT_E[0] & T725[0];
  assign T725[51] = ~T932[50];
  assign T725[50] = ~T932[49];
  assign T725[49] = ~T932[48];
  assign T725[48] = ~T932[47];
  assign T725[47] = ~T932[46];
  assign T725[46] = ~T932[45];
  assign T725[45] = ~T932[44];
  assign T725[44] = ~T932[43];
  assign T725[43] = ~T932[42];
  assign T725[42] = ~T932[41];
  assign T725[41] = ~T932[40];
  assign T725[40] = ~T932[39];
  assign T725[39] = ~T932[38];
  assign T725[38] = ~T932[37];
  assign T725[37] = ~T932[36];
  assign T725[36] = ~T932[35];
  assign T725[35] = ~T932[34];
  assign T725[34] = ~T932[33];
  assign T725[33] = ~T932[32];
  assign T725[32] = ~T932[31];
  assign T725[31] = ~T932[30];
  assign T725[30] = ~T932[29];
  assign T725[29] = ~T932[28];
  assign T725[28] = ~T932[27];
  assign T725[27] = ~T932[26];
  assign T725[26] = ~T932[25];
  assign T725[25] = ~T932[24];
  assign T725[24] = ~T932[23];
  assign T725[23] = ~T932[22];
  assign T725[22] = ~T932[21];
  assign T725[21] = ~T932[20];
  assign T725[20] = ~T932[19];
  assign T725[19] = ~T932[18];
  assign T725[18] = ~T932[17];
  assign T725[17] = ~T932[16];
  assign T725[16] = ~T932[15];
  assign T725[15] = ~T932[14];
  assign T725[14] = ~T932[13];
  assign T725[13] = ~T932[12];
  assign T725[12] = ~T932[11];
  assign T725[11] = ~T932[10];
  assign T725[10] = ~T932[9];
  assign T725[9] = ~T932[8];
  assign T725[8] = ~T932[7];
  assign T725[7] = ~T932[6];
  assign T725[6] = ~T932[5];
  assign T725[5] = ~T932[4];
  assign T725[4] = ~T586[0];
  assign T725[3] = ~T586[1];
  assign T725[2] = ~T586[2];
  assign T725[1] = ~T586[3];
  assign T725[0] = ~roundMask_E[0];
  assign N162 = ~sign_PC;
  assign T728[53] = sigAdjT_E[53] | 1'b0;
  assign T728[52] = sigAdjT_E[52] | T932[51];
  assign T728[51] = sigAdjT_E[51] | T932[50];
  assign T728[50] = sigAdjT_E[50] | T932[49];
  assign T728[49] = sigAdjT_E[49] | T932[48];
  assign T728[48] = sigAdjT_E[48] | T932[47];
  assign T728[47] = sigAdjT_E[47] | T932[46];
  assign T728[46] = sigAdjT_E[46] | T932[45];
  assign T728[45] = sigAdjT_E[45] | T932[44];
  assign T728[44] = sigAdjT_E[44] | T932[43];
  assign T728[43] = sigAdjT_E[43] | T932[42];
  assign T728[42] = sigAdjT_E[42] | T932[41];
  assign T728[41] = sigAdjT_E[41] | T932[40];
  assign T728[40] = sigAdjT_E[40] | T932[39];
  assign T728[39] = sigAdjT_E[39] | T932[38];
  assign T728[38] = sigAdjT_E[38] | T932[37];
  assign T728[37] = sigAdjT_E[37] | T932[36];
  assign T728[36] = sigAdjT_E[36] | T932[35];
  assign T728[35] = sigAdjT_E[35] | T932[34];
  assign T728[34] = sigAdjT_E[34] | T932[33];
  assign T728[33] = sigAdjT_E[33] | T932[32];
  assign T728[32] = sigAdjT_E[32] | T932[31];
  assign T728[31] = sigAdjT_E[31] | T932[30];
  assign T728[30] = sigAdjT_E[30] | T932[29];
  assign T728[29] = sigAdjT_E[29] | T932[28];
  assign T728[28] = sigAdjT_E[28] | T932[27];
  assign T728[27] = sigAdjT_E[27] | T932[26];
  assign T728[26] = sigAdjT_E[26] | T932[25];
  assign T728[25] = sigAdjT_E[25] | T932[24];
  assign T728[24] = sigAdjT_E[24] | T932[23];
  assign T728[23] = sigAdjT_E[23] | T932[22];
  assign T728[22] = sigAdjT_E[22] | T932[21];
  assign T728[21] = sigAdjT_E[21] | T932[20];
  assign T728[20] = sigAdjT_E[20] | T932[19];
  assign T728[19] = sigAdjT_E[19] | T932[18];
  assign T728[18] = sigAdjT_E[18] | T932[17];
  assign T728[17] = sigAdjT_E[17] | T932[16];
  assign T728[16] = sigAdjT_E[16] | T932[15];
  assign T728[15] = sigAdjT_E[15] | T932[14];
  assign T728[14] = sigAdjT_E[14] | T932[13];
  assign T728[13] = sigAdjT_E[13] | T932[12];
  assign T728[12] = sigAdjT_E[12] | T932[11];
  assign T728[11] = sigAdjT_E[11] | T932[10];
  assign T728[10] = sigAdjT_E[10] | T932[9];
  assign T728[9] = sigAdjT_E[9] | T932[8];
  assign T728[8] = sigAdjT_E[8] | T932[7];
  assign T728[7] = sigAdjT_E[7] | T932[6];
  assign T728[6] = sigAdjT_E[6] | T932[5];
  assign T728[5] = sigAdjT_E[5] | T932[4];
  assign T728[4] = sigAdjT_E[4] | T586[0];
  assign T728[3] = sigAdjT_E[3] | T586[1];
  assign T728[2] = sigAdjT_E[2] | T586[2];
  assign T728[1] = sigAdjT_E[1] | T586[3];
  assign T728[0] = sigAdjT_E[0] | roundMask_E[0];
  assign T730 = T742 | T731;
  assign T731 = N411 & T732;
  assign T732 = T736 | T733;
  assign T733 = T734 & N409;
  assign T734 = extraT_E & T735;
  assign T735 = ~trueLtX_E1;
  assign T736 = N463 | T737;
  assign T737 = T740 & T738;
  assign T738 = ~roundMask_E[0];
  assign T740 = extraT_E | T741;
  assign T741 = ~trueLtX_E1;
  assign T742 = T753 | T743;
  assign T743 = T944[0] & T744;
  assign T744 = T749 | T745;
  assign T745 = ~all1sHiRoundT_E;
  assign all1sHiRoundT_E = T746 & N409;
  assign T746 = T747 | N463;
  assign T747 = ~roundMask_E[0];
  assign T749 = T751 & T750;
  assign T750 = ~isZeroRemT_E;
  assign T751 = extraT_E & T752;
  assign T752 = ~trueLtX_E1;
  assign T753 = T754 & all1sHiRoundT_E;
  assign T754 = T756 & T755;
  assign T755 = ~trueLtX_E1;
  assign T756 = roundMagDown_PC & extraT_E;
  assign roundMagDown_PC = T758 & T757;
  assign T757 = ~N411;
  assign T758 = ~T944[0];
  assign T759[13] = T766[13] | T760[13];
  assign T759[12] = T766[12] | T760[12];
  assign T759[11] = T766[11] | T760[11];
  assign T759[10] = T766[10] | T760[10];
  assign T759[9] = T766[9] | T760[9];
  assign T759[8] = T766[8] | T760[8];
  assign T759[7] = T766[7] | T760[7];
  assign T759[6] = T766[6] | T760[6];
  assign T759[5] = T766[5] | T760[5];
  assign T759[4] = T766[4] | T760[4];
  assign T759[3] = T766[3] | T760[3];
  assign T759[2] = T766[2] | T760[2];
  assign T759[1] = T766[1] | T760[1];
  assign T759[0] = T766[0] | T760[0];
  assign N163 = ~T761;
  assign T761 = T763 & T762;
  assign T762 = ~E_E_div;
  assign T763 = sigY_E1_53 & T764;
  assign T764 = ~sqrtOp_PC;
  assign T766[13] = T772[13] | T767[13];
  assign T766[12] = T772[12] | T767[12];
  assign T766[11] = T772[11] | T767[11];
  assign T766[10] = T772[10] | T767[10];
  assign T766[9] = T772[9] | T767[9];
  assign T766[8] = T772[8] | T767[8];
  assign T766[7] = T772[7] | T767[7];
  assign T766[6] = T772[6] | T767[6];
  assign T766[5] = T772[5] | T767[5];
  assign T766[4] = T772[4] | T767[4];
  assign T766[3] = T772[3] | T767[3];
  assign T766[2] = T772[2] | T767[2];
  assign T766[1] = T772[1] | T767[1];
  assign T766[0] = T772[0] | T767[0];
  assign N164 = ~T768;
  assign T768 = T769 & E_E_div;
  assign T769 = sigY_E1_53 & T770;
  assign T770 = ~sqrtOp_PC;
  assign N165 = ~T773;
  assign T773 = ~sigY_E1_53;
  assign io_exceptionFlags[2] = normalCase_PC & overflowY_E1;
  assign overflowY_E1 = T778 & T776;
  assign T778 = ~sExpY_E1[13];
  assign io_exceptionFlags[3] = T781 & N533;
  assign T781 = T783 & T782;
  assign T782 = ~N536;
  assign T783 = T785 & T784;
  assign T784 = ~N539;
  assign T785 = ~sqrtOp_PC;
  assign io_exceptionFlags[4] = T798 | notSigNaN_invalid_PC;
  assign T786 = T792 | T787;
  assign T787 = isInfA_PC & isInfB_PC;
  assign isInfB_PC = N540 & T788;
  assign T788 = ~specialCodeB_PC[0];
  assign isInfA_PC = N539 & T790;
  assign T790 = ~specialCodeA_PC[0];
  assign T792 = N536 & N533;
  assign T793 = T794 & sign_PC;
  assign T794 = T796 & T795;
  assign T795 = ~N533;
  assign T796 = ~isNaNB_PC;
  assign isNaNB_PC = N540 & specialCodeB_PC[0];
  assign T798 = T800 | isSigNaNB_PC;
  assign isSigNaNB_PC = isNaNB_PC & T799;
  assign T799 = ~sigB_PC[51];
  assign T800 = T809 & isSigNaNA_PC;
  assign isSigNaNA_PC = isNaNA_PC & T801;
  assign T801 = ~fractA_51_PC;
  assign isNaNA_PC = N539 & specialCodeA_PC[0];
  assign T809 = ~sqrtOp_PC;
  assign io_out[51] = T816[51] | T812[51];
  assign io_out[50] = T816[50] | 1'b0;
  assign io_out[49] = T816[49] | 1'b0;
  assign io_out[48] = T816[48] | 1'b0;
  assign io_out[47] = T816[47] | 1'b0;
  assign io_out[46] = T816[46] | 1'b0;
  assign io_out[45] = T816[45] | 1'b0;
  assign io_out[44] = T816[44] | 1'b0;
  assign io_out[43] = T816[43] | 1'b0;
  assign io_out[42] = T816[42] | 1'b0;
  assign io_out[41] = T816[41] | 1'b0;
  assign io_out[40] = T816[40] | 1'b0;
  assign io_out[39] = T816[39] | 1'b0;
  assign io_out[38] = T816[38] | 1'b0;
  assign io_out[37] = T816[37] | 1'b0;
  assign io_out[36] = T816[36] | 1'b0;
  assign io_out[35] = T816[35] | 1'b0;
  assign io_out[34] = T816[34] | 1'b0;
  assign io_out[33] = T816[33] | 1'b0;
  assign io_out[32] = T816[32] | 1'b0;
  assign io_out[31] = T816[31] | 1'b0;
  assign io_out[30] = T816[30] | 1'b0;
  assign io_out[29] = T816[29] | 1'b0;
  assign io_out[28] = T816[28] | 1'b0;
  assign io_out[27] = T816[27] | 1'b0;
  assign io_out[26] = T816[26] | 1'b0;
  assign io_out[25] = T816[25] | 1'b0;
  assign io_out[24] = T816[24] | 1'b0;
  assign io_out[23] = T816[23] | 1'b0;
  assign io_out[22] = T816[22] | 1'b0;
  assign io_out[21] = T816[21] | 1'b0;
  assign io_out[20] = T816[20] | 1'b0;
  assign io_out[19] = T816[19] | 1'b0;
  assign io_out[18] = T816[18] | 1'b0;
  assign io_out[17] = T816[17] | 1'b0;
  assign io_out[16] = T816[16] | 1'b0;
  assign io_out[15] = T816[15] | 1'b0;
  assign io_out[14] = T816[14] | 1'b0;
  assign io_out[13] = T816[13] | 1'b0;
  assign io_out[12] = T816[12] | 1'b0;
  assign io_out[11] = T816[11] | 1'b0;
  assign io_out[10] = T816[10] | 1'b0;
  assign io_out[9] = T816[9] | 1'b0;
  assign io_out[8] = T816[8] | 1'b0;
  assign io_out[7] = T816[7] | 1'b0;
  assign io_out[6] = T816[6] | 1'b0;
  assign io_out[5] = T816[5] | 1'b0;
  assign io_out[4] = T816[4] | 1'b0;
  assign io_out[3] = T816[3] | 1'b0;
  assign io_out[2] = T816[2] | 1'b0;
  assign io_out[1] = T816[1] | 1'b0;
  assign io_out[0] = T816[0] | 1'b0;
  assign T812[51] = T813 | notSigNaN_invalid_PC;
  assign T813 = T814 | isNaNB_PC;
  assign T814 = T815 & isNaNA_PC;
  assign T815 = ~sqrtOp_PC;
  assign T816[51] = T819[51] | T817[51];
  assign T816[50] = T819[50] | T817[51];
  assign T816[49] = T819[49] | T817[51];
  assign T816[48] = T819[48] | T817[51];
  assign T816[47] = T819[47] | T817[51];
  assign T816[46] = T819[46] | T817[51];
  assign T816[45] = T819[45] | T817[51];
  assign T816[44] = T819[44] | T817[51];
  assign T816[43] = T819[43] | T817[51];
  assign T816[42] = T819[42] | T817[51];
  assign T816[41] = T819[41] | T817[51];
  assign T816[40] = T819[40] | T817[51];
  assign T816[39] = T819[39] | T817[51];
  assign T816[38] = T819[38] | T817[51];
  assign T816[37] = T819[37] | T817[51];
  assign T816[36] = T819[36] | T817[51];
  assign T816[35] = T819[35] | T817[51];
  assign T816[34] = T819[34] | T817[51];
  assign T816[33] = T819[33] | T817[51];
  assign T816[32] = T819[32] | T817[51];
  assign T816[31] = T819[31] | T817[51];
  assign T816[30] = T819[30] | T817[51];
  assign T816[29] = T819[29] | T817[51];
  assign T816[28] = T819[28] | T817[51];
  assign T816[27] = T819[27] | T817[51];
  assign T816[26] = T819[26] | T817[51];
  assign T816[25] = T819[25] | T817[51];
  assign T816[24] = T819[24] | T817[51];
  assign T816[23] = T819[23] | T817[51];
  assign T816[22] = T819[22] | T817[51];
  assign T816[21] = T819[21] | T817[51];
  assign T816[20] = T819[20] | T817[51];
  assign T816[19] = T819[19] | T817[51];
  assign T816[18] = T819[18] | T817[51];
  assign T816[17] = T819[17] | T817[51];
  assign T816[16] = T819[16] | T817[51];
  assign T816[15] = T819[15] | T817[51];
  assign T816[14] = T819[14] | T817[51];
  assign T816[13] = T819[13] | T817[51];
  assign T816[12] = T819[12] | T817[51];
  assign T816[11] = T819[11] | T817[51];
  assign T816[10] = T819[10] | T817[51];
  assign T816[9] = T819[9] | T817[51];
  assign T816[8] = T819[8] | T817[51];
  assign T816[7] = T819[7] | T817[51];
  assign T816[6] = T819[6] | T817[51];
  assign T816[5] = T819[5] | T817[51];
  assign T816[4] = T819[4] | T817[51];
  assign T816[3] = T819[3] | T817[51];
  assign T816[2] = T819[2] | T817[51];
  assign T816[1] = T819[1] | T817[51];
  assign T816[0] = T819[0] | T817_0;
  assign T946[0] = io_exceptionFlags[2] & T818;
  assign T818 = ~overflowY_roundMagUp_PC;
  assign overflowY_roundMagUp_PC = N411 | T944[0];
  assign N166 = ~T820;
  assign T820 = T821 | T812[51];
  assign T821 = notSpecial_isZeroOut_E1 | totalUnderflowY_E1;
  assign T822 = T825 | T823;
  assign T823 = totalUnderflowY_E1 & T824;
  assign T824 = ~T944[0];
  assign T825 = N536 | isInfB_PC;
  assign io_out[63] = T827[11] | T826[11];
  assign io_out[62] = T827[10] | T826[11];
  assign io_out[61] = T827[9] | T826[11];
  assign io_out[60] = T827[8] | 1'b0;
  assign io_out[59] = T827[7] | 1'b0;
  assign io_out[58] = T827[6] | 1'b0;
  assign io_out[57] = T827[5] | 1'b0;
  assign io_out[56] = T827[4] | 1'b0;
  assign io_out[55] = T827[3] | 1'b0;
  assign io_out[54] = T827[2] | 1'b0;
  assign io_out[53] = T827[1] | 1'b0;
  assign io_out[52] = T827[0] | 1'b0;
  assign T826[11] = T812[51];
  assign T827[11] = T832[11] | T828[11];
  assign T827[10] = T832[10] | T828[11];
  assign T827[9] = T832[9] | 1'b0;
  assign T827[8] = T832[8] | 1'b0;
  assign T827[7] = T832[7] | 1'b0;
  assign T827[6] = T832[6] | 1'b0;
  assign T827[5] = T832[5] | 1'b0;
  assign T827[4] = T832[4] | 1'b0;
  assign T827[3] = T832[3] | 1'b0;
  assign T827[2] = T832[2] | 1'b0;
  assign T827[1] = T832[1] | 1'b0;
  assign T827[0] = T832[0] | 1'b0;
  assign T828[11] = notNaN_isInfOut_E1;
  assign T829 = T831 | T830;
  assign T830 = io_exceptionFlags[2] & overflowY_roundMagUp_PC;
  assign T831 = isInfA_PC | N533;
  assign T832[11] = T834[11] | T833[11];
  assign T832[10] = T834[10] | 1'b0;
  assign T832[9] = T834[9] | T833[11];
  assign T832[8] = T834[8] | T833[11];
  assign T832[7] = T834[7] | T833[11];
  assign T832[6] = T834[6] | T833[11];
  assign T832[5] = T834[5] | T833[11];
  assign T832[4] = T834[4] | T833[11];
  assign T832[3] = T834[3] | T833[11];
  assign T832[2] = T834[2] | T833[11];
  assign T832[1] = T834[1] | T833[11];
  assign T832[0] = T834[0] | T833[11];
  assign T833[11] = T946[0];
  assign T834[11] = T837[11] | 1'b0;
  assign T834[10] = T837[10] | 1'b0;
  assign T834[9] = T837[9] | T835[9];
  assign T834[8] = T837[8] | T835[9];
  assign T834[7] = T837[7] | T835[9];
  assign T834[6] = T837[6] | T835[9];
  assign T834[5] = T837[5] | 1'b0;
  assign T834[4] = T837[4] | 1'b0;
  assign T834[3] = T837[3] | T835[9];
  assign T834[2] = T837[2] | T835[9];
  assign T834[1] = T837[1] | T835[9];
  assign T834[0] = T837[0] | 1'b0;
  assign T835[9] = pegMinFiniteMagOut_E1;
  assign pegMinFiniteMagOut_E1 = T836 & T944[0];
  assign T836 = normalCase_PC & totalUnderflowY_E1;
  assign T837[11] = T840[11] & T838[11];
  assign T837[10] = T840[10] & T838[10];
  assign T837[9] = T840[9] & T838[9];
  assign T837[8] = T840[8] & T838[8];
  assign T837[7] = T840[7] & T838[7];
  assign T837[6] = T840[6] & T838[6];
  assign T837[5] = T840[5] & T838[5];
  assign T837[4] = T840[4] & T838[4];
  assign T837[3] = T840[3] & T838[3];
  assign T837[2] = T840[2] & T838[2];
  assign T837[1] = T840[1] & T838[1];
  assign T837[0] = T840[0] & T838[0];
  assign T838[11] = ~1'b0;
  assign T838[10] = ~1'b0;
  assign T838[9] = ~T839[9];
  assign T838[8] = ~1'b0;
  assign T838[7] = ~1'b0;
  assign T838[6] = ~1'b0;
  assign T838[5] = ~1'b0;
  assign T838[4] = ~1'b0;
  assign T838[3] = ~1'b0;
  assign T838[2] = ~1'b0;
  assign T838[1] = ~1'b0;
  assign T838[0] = ~1'b0;
  assign T839[9] = notNaN_isInfOut_E1;
  assign T840[11] = T843[11] & T841[11];
  assign T840[10] = T843[10] & T841[10];
  assign T840[9] = T843[9] & T841[9];
  assign T840[8] = T843[8] & T841[8];
  assign T840[7] = T843[7] & T841[7];
  assign T840[6] = T843[6] & T841[6];
  assign T840[5] = T843[5] & T841[5];
  assign T840[4] = T843[4] & T841[4];
  assign T840[3] = T843[3] & T841[3];
  assign T840[2] = T843[2] & T841[2];
  assign T840[1] = T843[1] & T841[1];
  assign T840[0] = T843[0] & T841[0];
  assign T841[11] = ~1'b0;
  assign T841[10] = ~T842[10];
  assign T841[9] = ~1'b0;
  assign T841[8] = ~1'b0;
  assign T841[7] = ~1'b0;
  assign T841[6] = ~1'b0;
  assign T841[5] = ~1'b0;
  assign T841[4] = ~1'b0;
  assign T841[3] = ~1'b0;
  assign T841[2] = ~1'b0;
  assign T841[1] = ~1'b0;
  assign T841[0] = ~1'b0;
  assign T842[10] = T946[0];
  assign T843[11] = T846[11] & T844[11];
  assign T843[10] = T846[10] & T844[10];
  assign T843[9] = T846[9] & T844[9];
  assign T843[8] = T846[8] & T844[8];
  assign T843[7] = T846[7] & T844[7];
  assign T843[6] = T846[6] & T844[6];
  assign T843[5] = T846[5] & T844[5];
  assign T843[4] = T846[4] & T844[4];
  assign T843[3] = T846[3] & T844[3];
  assign T843[2] = T846[2] & T844[2];
  assign T843[1] = T846[1] & T844[1];
  assign T843[0] = T846[0] & T844[0];
  assign T844[11] = ~T845[11];
  assign T844[10] = ~T845[11];
  assign T844[9] = ~1'b0;
  assign T844[8] = ~1'b0;
  assign T844[7] = ~1'b0;
  assign T844[6] = ~1'b0;
  assign T844[5] = ~T845[11];
  assign T844[4] = ~T845[11];
  assign T844[3] = ~1'b0;
  assign T844[2] = ~1'b0;
  assign T844[1] = ~1'b0;
  assign T844[0] = ~T845[11];
  assign T845[11] = pegMinFiniteMagOut_E1;
  assign T846[11] = T709[11] & T847[11];
  assign T846[10] = T709[10] & T847[10];
  assign T846[9] = T709[9] & T847[9];
  assign T846[8] = T709[8] & T847[8];
  assign T846[7] = T709[7] & T847[7];
  assign T846[6] = T709[6] & T847[6];
  assign T846[5] = T709[5] & T847[5];
  assign T846[4] = T709[4] & T847[4];
  assign T846[3] = T709[3] & T847[3];
  assign T846[2] = T709[2] & T847[2];
  assign T846[1] = T709[1] & T847[1];
  assign T846[0] = T709[0] & T847[0];
  assign T847[11] = ~T848[11];
  assign T847[10] = ~T848[11];
  assign T847[9] = ~T848[11];
  assign T847[8] = ~1'b0;
  assign T847[7] = ~1'b0;
  assign T847[6] = ~1'b0;
  assign T847[5] = ~1'b0;
  assign T847[4] = ~1'b0;
  assign T847[3] = ~1'b0;
  assign T847[2] = ~1'b0;
  assign T847[1] = ~1'b0;
  assign T847[0] = ~1'b0;
  assign T848[11] = notSpecial_isZeroOut_E1;
  assign io_out[64] = T851 & T849;
  assign T850 = N533 & sign_PC;
  assign T851 = ~T812[51];
  assign io_outValid_sqrt = leaving_PC & sqrtOp_PC;
  assign io_outValid_div = leaving_PC & T854;
  assign T854 = ~sqrtOp_PC;
  assign io_inReady_sqrt = T857 & T856;
  assign T856 = ~cyc_B1_sqrt;
  assign T857 = T859 & T858;
  assign T858 = ~cyc_B2_div;
  assign T859 = T861 & T860;
  assign T860 = ~cyc_B4_sqrt;
  assign T861 = T863 & T862;
  assign T862 = ~cyc_B5_sqrt;
  assign T863 = ready_PA & T864;
  assign T864 = ~cyc_B6_sqrt;
  assign ready_PA = T866 | valid_leaving_PA;
  assign T866 = ~valid_PA;
  assign io_inReady_div = T869 & T868;
  assign T868 = ~N476;
  assign T869 = T871 & T870;
  assign T870 = ~N481;
  assign T871 = T873 & T872;
  assign T872 = ~cyc_B1_sqrt;
  assign T873 = T875 & T874;
  assign T874 = ~N485;
  assign T875 = T877 & T876;
  assign T876 = ~N493;
  assign T877 = T879 & T878;
  assign T878 = ~cyc_B4_sqrt;
  assign T879 = T881 & T880;
  assign T880 = ~cyc_B5_sqrt;
  assign T881 = T883 & T882;
  assign T882 = ~cyc_B6_sqrt;
  assign T883 = ready_PA & T884;
  assign T884 = ~N506;
  assign N167 = T30 | reset;
  assign N168 = ~N167;
  assign N173 = T67 | reset;
  assign N174 = ~N173;
  assign N177 = T106 | reset;
  assign N178 = ~N177;
  assign N183 = T104 | reset;
  assign N184 = ~N183;
  assign N190 = T102 | reset;
  assign N191 = ~N190;
  assign N196 = T124 | reset;
  assign N197 = ~N196;
  assign N200 = T155 | reset;
  assign N201 = ~N200;
  assign N204 = ~reset;
  assign N205 = T30 & N204;
  assign N206 = T67 & N204;
  assign N207 = T106 & N204;
  assign N208 = T104 & N204;
  assign N209 = T102 & N204;
  assign N210 = T124 & N204;
  assign N211 = T155 & N204;
  assign N212 = ~N323;

endmodule