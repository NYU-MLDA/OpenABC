module csr_regfile_0000000000000000_1
(
  clk_i,
  rst_ni,
  time_irq_i,
  flush_o,
  halt_csr_o,
  commit_instr_i,
  commit_ack_i,
  boot_addr_i,
  hart_id_i,
  ex_i,
  csr_op_i,
  csr_addr_i,
  csr_wdata_i,
  csr_rdata_o,
  dirty_fp_state_i,
  csr_write_fflags_i,
  pc_i,
  csr_exception_o,
  epc_o,
  eret_o,
  trap_vector_base_o,
  priv_lvl_o,
  fs_o,
  fflags_o,
  frm_o,
  fprec_o,
  en_translation_o,
  en_ld_st_translation_o,
  ld_st_priv_lvl_o,
  sum_o,
  mxr_o,
  satp_ppn_o,
  asid_o,
  irq_i,
  ipi_i,
  debug_req_i,
  set_debug_pc_o,
  tvm_o,
  tw_o,
  tsr_o,
  debug_mode_o,
  single_step_o,
  icache_en_o,
  dcache_en_o,
  perf_addr_o,
  perf_data_o,
  perf_data_i,
  perf_we_o
);

  input [723:0] commit_instr_i;
  input [1:0] commit_ack_i;
  input [63:0] boot_addr_i;
  input [63:0] hart_id_i;
  input [128:0] ex_i;
  input [6:0] csr_op_i;
  input [11:0] csr_addr_i;
  input [63:0] csr_wdata_i;
  output [63:0] csr_rdata_o;
  input [63:0] pc_i;
  output [128:0] csr_exception_o;
  output [63:0] epc_o;
  output [63:0] trap_vector_base_o;
  output [1:0] priv_lvl_o;
  output [1:0] fs_o;
  output [4:0] fflags_o;
  output [2:0] frm_o;
  output [6:0] fprec_o;
  output [1:0] ld_st_priv_lvl_o;
  output [43:0] satp_ppn_o;
  output [0:0] asid_o;
  input [1:0] irq_i;
  output [4:0] perf_addr_o;
  output [63:0] perf_data_o;
  input [63:0] perf_data_i;
  input clk_i;
  input rst_ni;
  input time_irq_i;
  input dirty_fp_state_i;
  input csr_write_fflags_i;
  input ipi_i;
  input debug_req_i;
  output flush_o;
  output halt_csr_o;
  output eret_o;
  output en_translation_o;
  output en_ld_st_translation_o;
  output sum_o;
  output mxr_o;
  output set_debug_pc_o;
  output tvm_o;
  output tw_o;
  output tsr_o;
  output debug_mode_o;
  output single_step_o;
  output icache_en_o;
  output dcache_en_o;
  output perf_we_o;
  wire [63:0] csr_rdata_o,epc_o,trap_vector_base_o,perf_data_o,csr_wdata,cycle_d,dpc_d,
  dscratch0_d,dscratch1_d,mtvec_d,mie_d,mepc_d,mcause_d,mscratch_d,mtval_d,dcache_d,
  icache_d,sepc_d,scause_d,stvec_d,sscratch_d,stval_d,satp_d;
  wire [128:0] csr_exception_o;
  wire [1:0] priv_lvl_o,ld_st_priv_lvl_o,priv_lvl_d;
  wire [4:0] perf_addr_o;
  wire flush_o,eret_o,en_translation_o,set_debug_pc_o,icache_en_o,perf_we_o,N0,N1,N2,
  N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,
  N168,csr_read,read_access_exception,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,
  N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,
  N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,
  N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
  N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,
  N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,
  N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,
  N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
  N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,
  N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,
  N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,
  N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,
  N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,
  N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,
  N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,
  N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,
  N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,
  N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,
  N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
  N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
  N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,
  N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,
  N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,
  N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,
  N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,
  N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,
  N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,
  N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,
  N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
  N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,
  N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,
  N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,
  N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,
  N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,
  N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,
  N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,
  N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,
  N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,
  N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,
  N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,
  N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,
  N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,
  N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,
  N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,
  N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,csr_we,mprv,mret,
  sret,dret,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,
  N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,
  N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,
  N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,
  N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,
  N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,
  N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,
  N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,
  N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,
  N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,
  N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,
  N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,
  N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,
  N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,
  N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,
  N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,
  N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,
  N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,
  N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,
  N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,
  N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,
  N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,
  N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,
  N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,
  N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,
  N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,
  N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,
  N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,
  N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,
  N1417,N1418,N1419,N1420,update_access_exception,fcsr_d_fprec__6_,
  fcsr_d_fprec__5_,fcsr_d_fprec__4_,fcsr_d_fprec__3_,fcsr_d_fprec__2_,fcsr_d_fprec__1_,
  fcsr_d_fprec__0_,fcsr_d_frm__2_,fcsr_d_frm__1_,fcsr_d_frm__0_,fcsr_d_fflags__4_,
  fcsr_d_fflags__3_,fcsr_d_fflags__2_,fcsr_d_fflags__1_,fcsr_d_fflags__0_,debug_mode_d,
  mstatus_d_sd_,mstatus_d_wpri4__62_,mstatus_d_wpri4__61_,mstatus_d_wpri4__60_,
  mstatus_d_wpri4__59_,mstatus_d_wpri4__58_,mstatus_d_wpri4__57_,mstatus_d_wpri4__56_,
  mstatus_d_wpri4__55_,mstatus_d_wpri4__54_,mstatus_d_wpri4__53_,mstatus_d_wpri4__52_,
  mstatus_d_wpri4__51_,mstatus_d_wpri4__50_,mstatus_d_wpri4__49_,
  mstatus_d_wpri4__48_,mstatus_d_wpri4__47_,mstatus_d_wpri4__46_,mstatus_d_wpri4__45_,
  mstatus_d_wpri4__44_,mstatus_d_wpri4__43_,mstatus_d_wpri4__42_,mstatus_d_wpri4__41_,
  mstatus_d_wpri4__40_,mstatus_d_wpri4__39_,mstatus_d_wpri4__38_,mstatus_d_wpri4__37_,
  mstatus_d_wpri4__36_,mstatus_d_wpri3__8_,mstatus_d_wpri3__7_,mstatus_d_wpri3__6_,
  mstatus_d_wpri3__5_,mstatus_d_wpri3__4_,mstatus_d_wpri3__3_,mstatus_d_wpri3__2_,
  mstatus_d_wpri3__1_,mstatus_d_wpri3__0_,mstatus_d_tsr_,mstatus_d_tw_,mstatus_d_tvm_,
  mstatus_d_mxr_,mstatus_d_sum_,mstatus_d_mprv_,mstatus_d_xs__1_,mstatus_d_xs__0_,
  mstatus_d_fs__1_,mstatus_d_fs__0_,mstatus_d_mpp__1_,mstatus_d_mpp__0_,
  mstatus_d_wpri2__1_,mstatus_d_wpri2__0_,mstatus_d_spp_,mstatus_d_mpie_,mstatus_d_wpri1_,
  mstatus_d_spie_,mstatus_d_upie_,mstatus_d_mie_,mstatus_d_wpri0_,mstatus_d_sie_,
  mstatus_d_uie_,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,
  N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,
  N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,
  N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,
  N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,
  N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,
  N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,mip_d_9,
  mip_d_5,mip_d_1,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,
  N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
  N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,
  N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,
  N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,
  N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,
  N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,
  N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,
  N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,
  N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,
  N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,
  N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,
  N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,
  N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,
  N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,
  N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,
  N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,
  N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,
  N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,
  N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,
  N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,
  N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,
  N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,
  N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
  N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,
  N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,
  N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,
  N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,
  N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,
  N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,
  N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
  N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,
  N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,
  N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,
  N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,
  N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,
  N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,
  N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,
  N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,
  N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,
  N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,
  N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,
  N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,
  N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,
  N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,
  N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,
  N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,
  N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,
  N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,
  N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,
  N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
  N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,
  N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,
  N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,
  N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,
  N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,
  N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,
  N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,
  N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,
  N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,
  N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,
  N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,
  N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,
  N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,
  N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,
  N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,
  N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,
  N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,
  N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,
  N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,
  N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,
  N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,
  N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,
  N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,
  N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,
  N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,
  N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,
  N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,
  N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,
  N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,
  N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,
  N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,
  N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,
  N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,
  N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,
  N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,
  N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,
  N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,
  N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,
  N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,
  N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,
  N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,
  N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,
  N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,
  N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,
  N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,
  N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,
  N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,
  N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,
  N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,
  N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,
  N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,
  N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,
  N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,
  N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,
  N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,
  N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,
  N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
  N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,
  N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,
  N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,
  N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,
  N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,
  N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,
  N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,
  N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,
  N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,
  N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,
  N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,
  N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,
  N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,
  N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,
  N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,
  N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,
  N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,
  N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,
  N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,
  N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,
  N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,
  N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,
  N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,
  N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,
  N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,
  N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,
  N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,
  N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,
  N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,
  N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,
  N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,
  N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,
  N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,
  N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,
  N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,
  N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,
  N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,
  N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,
  N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,
  N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,
  N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,
  N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,
  N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,
  N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,
  N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,
  N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,
  N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,
  N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,
  N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,
  N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,
  N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,
  N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,
  N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,
  N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,
  N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,
  N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,
  N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,
  N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,
  N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,
  N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,
  N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,
  N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,
  N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,
  N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,
  N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,
  N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,
  N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,
  N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,
  N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,
  N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,
  N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,
  N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,
  N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,
  N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,
  N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,
  N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,
  N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,
  N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,
  N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
  N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,
  N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,
  N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,
  N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,
  N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,
  N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,
  N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,
  N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,
  N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,
  N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,
  N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,
  N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,
  N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,
  N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,
  N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,
  N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,
  N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,
  N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,
  N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,
  N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,
  N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,
  N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,
  N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,
  N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,
  N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,
  N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,
  N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,
  N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,
  N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,
  N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,
  N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,
  N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,
  N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,
  N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
  N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,
  N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,
  N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,
  N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,N4558,N4559,N4560,
  N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,
  N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,
  N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,N4598,N4599,N4600,
  N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,
  N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,
  N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,
  N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,
  N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,
  N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4680,
  N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,
  N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,
  N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718,N4719,N4720,
  N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,
  N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,
  N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,
  N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,
  N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,
  N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,N4798,N4799,N4800,
  N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,
  N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,
  N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,N4838,N4839,N4840,
  N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,
  N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,
  N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,N4878,N4879,N4880,
  N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,
  N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,
  N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920,
  N4921,en_ld_st_translation_d,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,N4930,
  N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,
  N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,
  N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,N4970,
  N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,
  N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,
  N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,N5010,
  N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,
  N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,
  N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,N5050,
  N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,
  N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,
  N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,
  N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,
  N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,
  N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,
  N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,
  N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,
  N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,N5170,
  N5171,wfi_d,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,
  N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,
  N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,
  N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,
  N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,
  N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,
  N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,
  N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,
  N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,
  N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,
  N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,
  N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,
  N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,
  N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,
  N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,
  N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,
  N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,
  N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,
  N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,
  N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,
  N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,
  N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,
  N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,
  N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,
  N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,
  N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,
  N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,
  N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,
  N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,
  N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,
  N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,
  N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,
  N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,
  N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,
  N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,
  N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,
  N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,
  N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,
  N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,
  N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,
  N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,
  N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,
  N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,
  N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,
  N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,
  N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,
  N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,
  N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,
  N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,
  N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,
  N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,
  N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,
  N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,
  N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,
  N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,
  N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,
  N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,
  N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,
  N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,
  N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,
  N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,
  N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,
  N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,
  N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,
  N6023,N6024,N6025,N6026,N6027,N6028;
  wire [9:9] csr_rdata;
  wire [31:0] dcsr_d;
  wire [1:1] trap_to_priv_lvl;
  reg halt_csr_o,debug_mode_o,dcsr_q_xdebugver__31_,dcsr_q_xdebugver__30_,
  dcsr_q_xdebugver__29_,dcsr_q_xdebugver__28_,dcsr_q_zero2__27_,dcsr_q_zero2__26_,
  dcsr_q_zero2__25_,dcsr_q_zero2__24_,dcsr_q_zero2__23_,dcsr_q_zero2__22_,dcsr_q_zero2__21_,
  dcsr_q_zero2__20_,dcsr_q_zero2__19_,dcsr_q_zero2__18_,dcsr_q_zero2__17_,
  dcsr_q_zero2__16_,dcsr_q_ebreakm_,dcsr_q_zero1_,dcsr_q_ebreaks_,dcsr_q_ebreaku_,
  dcsr_q_stepie_,dcsr_q_stopcount_,dcsr_q_stoptime_,dcsr_q_cause__8_,dcsr_q_cause__7_,
  dcsr_q_cause__6_,dcsr_q_zero0_,dcsr_q_mprven_,dcsr_q_nmip_,single_step_o,
  dcsr_q_prv__1_,dcsr_q_prv__0_,mstatus_q_sd_,mstatus_q_wpri4__62_,mstatus_q_wpri4__61_,
  mstatus_q_wpri4__60_,mstatus_q_wpri4__59_,mstatus_q_wpri4__58_,mstatus_q_wpri4__57_,
  mstatus_q_wpri4__56_,mstatus_q_wpri4__55_,mstatus_q_wpri4__54_,
  mstatus_q_wpri4__53_,mstatus_q_wpri4__52_,mstatus_q_wpri4__51_,mstatus_q_wpri4__50_,
  mstatus_q_wpri4__49_,mstatus_q_wpri4__48_,mstatus_q_wpri4__47_,mstatus_q_wpri4__46_,
  mstatus_q_wpri4__45_,mstatus_q_wpri4__44_,mstatus_q_wpri4__43_,mstatus_q_wpri4__42_,
  mstatus_q_wpri4__41_,mstatus_q_wpri4__40_,mstatus_q_wpri4__39_,mstatus_q_wpri4__38_,
  mstatus_q_wpri4__37_,mstatus_q_wpri4__36_,mstatus_q_sxl__1_,mstatus_q_sxl__0_,
  mstatus_q_uxl__1_,mstatus_q_uxl__0_,mstatus_q_wpri3__8_,mstatus_q_wpri3__7_,
  mstatus_q_wpri3__6_,mstatus_q_wpri3__5_,mstatus_q_wpri3__4_,mstatus_q_wpri3__3_,
  mstatus_q_wpri3__2_,mstatus_q_wpri3__1_,mstatus_q_wpri3__0_,tsr_o,tw_o,tvm_o,mxr_o,sum_o,
  mstatus_q_mprv_,mstatus_q_xs__1_,mstatus_q_xs__0_,mstatus_q_mpp__1_,
  mstatus_q_mpp__0_,mstatus_q_wpri2__1_,mstatus_q_wpri2__0_,mstatus_q_spp_,mstatus_q_mpie_,
  mstatus_q_wpri1_,mstatus_q_spie_,mstatus_q_upie_,mstatus_q_mie_,mstatus_q_wpri0_,
  mstatus_q_sie_,mstatus_q_uie_,mtvec_rst_load_q,medeleg_q_15,medeleg_q_8,
  medeleg_q_3,medeleg_q_0,mideleg_q_5,mideleg_q_1,mip_d_10,mip_q_9,mip_d_8,mip_q_7,mip_d_6,
  mip_q_5,mip_d_4,mip_q_3,mip_d_2,mip_q_1,mip_d_0,dcache_en_o,satp_q_mode__3_,
  satp_q_mode__2_,satp_q_mode__1_,satp_q_mode__0_,satp_q_asid__15_,satp_q_asid__14_,
  satp_q_asid__13_,satp_q_asid__12_,satp_q_asid__11_,satp_q_asid__10_,satp_q_asid__9_,
  satp_q_asid__8_,satp_q_asid__7_,satp_q_asid__6_,satp_q_asid__5_,satp_q_asid__4_,
  satp_q_asid__3_,satp_q_asid__2_,satp_q_asid__1_,en_ld_st_translation_o;
  reg [1:0] priv_lvl_q,fs_o;
  reg [6:0] fprec_o;
  reg [2:0] frm_o;
  reg [4:0] fflags_o;
  reg [63:0] dpc_q,dscratch0_q,dscratch1_q,mtvec_q,medeleg_d,mideleg_d,mie_q,mepc_q,mcause_q,
  mscratch_q,mtval_q,icache_q,sepc_q,scause_q,stvec_q,sscratch_q,stval_q,cycle_q,
  instret_q;
  reg [13:12] medeleg_q;
  reg [9:9] mideleg_q;
  reg [63:12] mip_d;
  reg [11:11] mip_q;
  reg [63:1] dcache_q;
  reg [0:0] asid_o;
  reg [43:0] satp_ppn_o;
  assign trap_vector_base_o[0] = 1'b0;
  assign trap_vector_base_o[1] = 1'b0;
  assign csr_exception_o[1] = 1'b0;
  assign csr_exception_o[2] = 1'b0;
  assign csr_exception_o[3] = 1'b0;
  assign csr_exception_o[4] = 1'b0;
  assign csr_exception_o[5] = 1'b0;
  assign csr_exception_o[6] = 1'b0;
  assign csr_exception_o[7] = 1'b0;
  assign csr_exception_o[8] = 1'b0;
  assign csr_exception_o[9] = 1'b0;
  assign csr_exception_o[10] = 1'b0;
  assign csr_exception_o[11] = 1'b0;
  assign csr_exception_o[12] = 1'b0;
  assign csr_exception_o[13] = 1'b0;
  assign csr_exception_o[14] = 1'b0;
  assign csr_exception_o[15] = 1'b0;
  assign csr_exception_o[16] = 1'b0;
  assign csr_exception_o[17] = 1'b0;
  assign csr_exception_o[18] = 1'b0;
  assign csr_exception_o[19] = 1'b0;
  assign csr_exception_o[20] = 1'b0;
  assign csr_exception_o[21] = 1'b0;
  assign csr_exception_o[22] = 1'b0;
  assign csr_exception_o[23] = 1'b0;
  assign csr_exception_o[24] = 1'b0;
  assign csr_exception_o[25] = 1'b0;
  assign csr_exception_o[26] = 1'b0;
  assign csr_exception_o[27] = 1'b0;
  assign csr_exception_o[28] = 1'b0;
  assign csr_exception_o[29] = 1'b0;
  assign csr_exception_o[30] = 1'b0;
  assign csr_exception_o[31] = 1'b0;
  assign csr_exception_o[32] = 1'b0;
  assign csr_exception_o[33] = 1'b0;
  assign csr_exception_o[34] = 1'b0;
  assign csr_exception_o[35] = 1'b0;
  assign csr_exception_o[36] = 1'b0;
  assign csr_exception_o[37] = 1'b0;
  assign csr_exception_o[38] = 1'b0;
  assign csr_exception_o[39] = 1'b0;
  assign csr_exception_o[40] = 1'b0;
  assign csr_exception_o[41] = 1'b0;
  assign csr_exception_o[42] = 1'b0;
  assign csr_exception_o[43] = 1'b0;
  assign csr_exception_o[44] = 1'b0;
  assign csr_exception_o[45] = 1'b0;
  assign csr_exception_o[46] = 1'b0;
  assign csr_exception_o[47] = 1'b0;
  assign csr_exception_o[48] = 1'b0;
  assign csr_exception_o[49] = 1'b0;
  assign csr_exception_o[50] = 1'b0;
  assign csr_exception_o[51] = 1'b0;
  assign csr_exception_o[52] = 1'b0;
  assign csr_exception_o[53] = 1'b0;
  assign csr_exception_o[54] = 1'b0;
  assign csr_exception_o[55] = 1'b0;
  assign csr_exception_o[56] = 1'b0;
  assign csr_exception_o[57] = 1'b0;
  assign csr_exception_o[58] = 1'b0;
  assign csr_exception_o[59] = 1'b0;
  assign csr_exception_o[60] = 1'b0;
  assign csr_exception_o[61] = 1'b0;
  assign csr_exception_o[62] = 1'b0;
  assign csr_exception_o[63] = 1'b0;
  assign csr_exception_o[64] = 1'b0;
  assign csr_exception_o[69] = 1'b0;
  assign csr_exception_o[70] = 1'b0;
  assign csr_exception_o[71] = 1'b0;
  assign csr_exception_o[72] = 1'b0;
  assign csr_exception_o[73] = 1'b0;
  assign csr_exception_o[74] = 1'b0;
  assign csr_exception_o[75] = 1'b0;
  assign csr_exception_o[76] = 1'b0;
  assign csr_exception_o[77] = 1'b0;
  assign csr_exception_o[78] = 1'b0;
  assign csr_exception_o[79] = 1'b0;
  assign csr_exception_o[80] = 1'b0;
  assign csr_exception_o[81] = 1'b0;
  assign csr_exception_o[82] = 1'b0;
  assign csr_exception_o[83] = 1'b0;
  assign csr_exception_o[84] = 1'b0;
  assign csr_exception_o[85] = 1'b0;
  assign csr_exception_o[86] = 1'b0;
  assign csr_exception_o[87] = 1'b0;
  assign csr_exception_o[88] = 1'b0;
  assign csr_exception_o[89] = 1'b0;
  assign csr_exception_o[90] = 1'b0;
  assign csr_exception_o[91] = 1'b0;
  assign csr_exception_o[92] = 1'b0;
  assign csr_exception_o[93] = 1'b0;
  assign csr_exception_o[94] = 1'b0;
  assign csr_exception_o[95] = 1'b0;
  assign csr_exception_o[96] = 1'b0;
  assign csr_exception_o[97] = 1'b0;
  assign csr_exception_o[98] = 1'b0;
  assign csr_exception_o[99] = 1'b0;
  assign csr_exception_o[100] = 1'b0;
  assign csr_exception_o[101] = 1'b0;
  assign csr_exception_o[102] = 1'b0;
  assign csr_exception_o[103] = 1'b0;
  assign csr_exception_o[104] = 1'b0;
  assign csr_exception_o[105] = 1'b0;
  assign csr_exception_o[106] = 1'b0;
  assign csr_exception_o[107] = 1'b0;
  assign csr_exception_o[108] = 1'b0;
  assign csr_exception_o[109] = 1'b0;
  assign csr_exception_o[110] = 1'b0;
  assign csr_exception_o[111] = 1'b0;
  assign csr_exception_o[112] = 1'b0;
  assign csr_exception_o[113] = 1'b0;
  assign csr_exception_o[114] = 1'b0;
  assign csr_exception_o[115] = 1'b0;
  assign csr_exception_o[116] = 1'b0;
  assign csr_exception_o[117] = 1'b0;
  assign csr_exception_o[118] = 1'b0;
  assign csr_exception_o[119] = 1'b0;
  assign csr_exception_o[120] = 1'b0;
  assign csr_exception_o[121] = 1'b0;
  assign csr_exception_o[122] = 1'b0;
  assign csr_exception_o[123] = 1'b0;
  assign csr_exception_o[124] = 1'b0;
  assign csr_exception_o[125] = 1'b0;
  assign csr_exception_o[126] = 1'b0;
  assign csr_exception_o[127] = 1'b0;
  assign perf_addr_o[4] = csr_addr_i[4];
  assign perf_addr_o[3] = csr_addr_i[3];
  assign perf_addr_o[2] = csr_addr_i[2];
  assign perf_addr_o[1] = csr_addr_i[1];
  assign perf_addr_o[0] = csr_addr_i[0];
  assign N171 = csr_addr_i[5] | csr_addr_i[4];
  assign N172 = csr_addr_i[3] | csr_addr_i[2];
  assign N173 = csr_addr_i[1] | N170;
  assign N174 = N5417 | N1859;
  assign N175 = N1860 | N171;
  assign N176 = N172 | N173;
  assign N177 = N174 | N175;
  assign N178 = N177 | N176;
  assign N181 = csr_addr_i[5] | csr_addr_i[4];
  assign N182 = csr_addr_i[3] | csr_addr_i[2];
  assign N183 = N180 | csr_addr_i[0];
  assign N184 = N1860 | N181;
  assign N185 = N182 | N183;
  assign N186 = N174 | N184;
  assign N187 = N186 | N185;
  assign N189 = csr_addr_i[5] | csr_addr_i[4];
  assign N190 = csr_addr_i[3] | csr_addr_i[2];
  assign N191 = N180 | N170;
  assign N192 = N1860 | N189;
  assign N193 = N190 | N191;
  assign N194 = N174 | N192;
  assign N195 = N194 | N193;
  assign N197 = N1857 | csr_addr_i[10];
  assign N198 = csr_addr_i[5] | csr_addr_i[4];
  assign N199 = csr_addr_i[3] | csr_addr_i[2];
  assign N200 = csr_addr_i[1] | csr_addr_i[0];
  assign N201 = N197 | N1859;
  assign N202 = N1860 | N198;
  assign N203 = N199 | N200;
  assign N204 = N201 | N202;
  assign N205 = N204 | N203;
  assign N207 = N5551 | csr_addr_i[6];
  assign N208 = N5552 | N5553;
  assign N209 = csr_addr_i[3] | csr_addr_i[2];
  assign N210 = csr_addr_i[1] | csr_addr_i[0];
  assign N211 = N207 | N208;
  assign N212 = N209 | N210;
  assign N213 = N1851 | N211;
  assign N214 = N213 | N212;
  assign N216 = N5552 | N5553;
  assign N217 = csr_addr_i[3] | csr_addr_i[2];
  assign N218 = csr_addr_i[1] | N170;
  assign N219 = N207 | N216;
  assign N220 = N217 | N218;
  assign N221 = N1851 | N219;
  assign N222 = N221 | N220;
  assign N224 = N5552 | N5553;
  assign N225 = csr_addr_i[3] | csr_addr_i[2];
  assign N226 = N180 | csr_addr_i[0];
  assign N227 = N207 | N224;
  assign N228 = N225 | N226;
  assign N229 = N1851 | N227;
  assign N230 = N229 | N228;
  assign N232 = N5552 | N5553;
  assign N233 = csr_addr_i[3] | csr_addr_i[2];
  assign N234 = N180 | N170;
  assign N235 = N207 | N232;
  assign N236 = N233 | N234;
  assign N237 = N1851 | N235;
  assign N238 = N237 | N236;
  assign N240 = N5552 | csr_addr_i[4];
  assign N241 = csr_addr_i[3] | csr_addr_i[2];
  assign N242 = csr_addr_i[1] | csr_addr_i[0];
  assign N243 = N207 | N240;
  assign N244 = N241 | N242;
  assign N245 = N1851 | N243;
  assign N246 = N245 | N244;
  assign N248 = N5552 | csr_addr_i[4];
  assign N249 = csr_addr_i[3] | csr_addr_i[2];
  assign N250 = csr_addr_i[1] | N170;
  assign N251 = N207 | N248;
  assign N252 = N249 | N250;
  assign N253 = N1851 | N251;
  assign N254 = N253 | N252;
  assign N256 = N5552 | csr_addr_i[4];
  assign N257 = csr_addr_i[3] | csr_addr_i[2];
  assign N258 = N180 | csr_addr_i[0];
  assign N259 = N207 | N256;
  assign N260 = N257 | N258;
  assign N261 = N1851 | N259;
  assign N262 = N261 | N260;
  assign N264 = N5552 | csr_addr_i[4];
  assign N265 = csr_addr_i[3] | csr_addr_i[2];
  assign N266 = N180 | N170;
  assign N267 = N207 | N264;
  assign N268 = N265 | N266;
  assign N269 = N1851 | N267;
  assign N270 = N269 | N268;
  assign N272 = csr_addr_i[5] | csr_addr_i[4];
  assign N273 = csr_addr_i[3] | csr_addr_i[2];
  assign N274 = csr_addr_i[1] | csr_addr_i[0];
  assign N275 = N1860 | N272;
  assign N276 = N273 | N274;
  assign N277 = N5423 | N275;
  assign N278 = N277 | N276;
  assign N281 = csr_addr_i[5] | csr_addr_i[4];
  assign N282 = csr_addr_i[3] | N280;
  assign N283 = csr_addr_i[1] | csr_addr_i[0];
  assign N284 = N1860 | N281;
  assign N285 = N282 | N283;
  assign N286 = N5423 | N284;
  assign N287 = N286 | N285;
  assign N289 = csr_addr_i[5] | csr_addr_i[4];
  assign N290 = csr_addr_i[3] | N280;
  assign N291 = csr_addr_i[1] | csr_addr_i[0];
  assign N292 = N5419 | N289;
  assign N293 = N290 | N291;
  assign N294 = N5423 | N292;
  assign N295 = N294 | N293;
  assign N297 = csr_addr_i[5] | csr_addr_i[4];
  assign N298 = csr_addr_i[3] | N280;
  assign N299 = csr_addr_i[1] | N170;
  assign N300 = N1860 | N297;
  assign N301 = N298 | N299;
  assign N302 = N5423 | N300;
  assign N303 = N302 | N301;
  assign N305 = csr_addr_i[5] | csr_addr_i[4];
  assign N306 = csr_addr_i[3] | N280;
  assign N307 = N180 | csr_addr_i[0];
  assign N308 = N1860 | N305;
  assign N309 = N306 | N307;
  assign N310 = N5423 | N308;
  assign N311 = N310 | N309;
  assign N313 = csr_addr_i[5] | csr_addr_i[4];
  assign N314 = csr_addr_i[3] | csr_addr_i[2];
  assign N315 = csr_addr_i[1] | csr_addr_i[0];
  assign N316 = N5419 | N313;
  assign N317 = N314 | N315;
  assign N318 = N5423 | N316;
  assign N319 = N318 | N317;
  assign N321 = csr_addr_i[5] | csr_addr_i[4];
  assign N322 = csr_addr_i[3] | csr_addr_i[2];
  assign N323 = csr_addr_i[1] | N170;
  assign N324 = N5419 | N321;
  assign N325 = N322 | N323;
  assign N326 = N5423 | N324;
  assign N327 = N326 | N325;
  assign N329 = csr_addr_i[5] | csr_addr_i[4];
  assign N330 = csr_addr_i[3] | csr_addr_i[2];
  assign N331 = N180 | csr_addr_i[0];
  assign N332 = N5419 | N329;
  assign N333 = N330 | N331;
  assign N334 = N5423 | N332;
  assign N335 = N334 | N333;
  assign N337 = csr_addr_i[5] | csr_addr_i[4];
  assign N338 = csr_addr_i[3] | csr_addr_i[2];
  assign N339 = N180 | N170;
  assign N340 = N5419 | N337;
  assign N341 = N338 | N339;
  assign N342 = N5423 | N340;
  assign N343 = N342 | N341;
  assign N345 = csr_addr_i[5] | csr_addr_i[4];
  assign N346 = csr_addr_i[3] | csr_addr_i[2];
  assign N347 = csr_addr_i[1] | csr_addr_i[0];
  assign N348 = N207 | N345;
  assign N349 = N346 | N347;
  assign N350 = N5423 | N348;
  assign N351 = N350 | N349;
  assign N353 = csr_addr_i[5] | csr_addr_i[4];
  assign N354 = csr_addr_i[3] | csr_addr_i[2];
  assign N355 = csr_addr_i[1] | csr_addr_i[0];
  assign N356 = N1860 | N353;
  assign N357 = N354 | N355;
  assign N358 = N5410 | N356;
  assign N359 = N358 | N357;
  assign N361 = csr_addr_i[5] | csr_addr_i[4];
  assign N362 = csr_addr_i[3] | csr_addr_i[2];
  assign N363 = csr_addr_i[1] | N170;
  assign N364 = N1860 | N361;
  assign N365 = N362 | N363;
  assign N366 = N5410 | N364;
  assign N367 = N366 | N365;
  assign N369 = csr_addr_i[5] | csr_addr_i[4];
  assign N370 = csr_addr_i[3] | csr_addr_i[2];
  assign N371 = N180 | csr_addr_i[0];
  assign N372 = N1860 | N369;
  assign N373 = N370 | N371;
  assign N374 = N5410 | N372;
  assign N375 = N374 | N373;
  assign N377 = csr_addr_i[5] | csr_addr_i[4];
  assign N378 = csr_addr_i[3] | csr_addr_i[2];
  assign N379 = N180 | N170;
  assign N380 = N1860 | N377;
  assign N381 = N378 | N379;
  assign N382 = N5410 | N380;
  assign N383 = N382 | N381;
  assign N385 = csr_addr_i[5] | csr_addr_i[4];
  assign N386 = csr_addr_i[3] | N280;
  assign N387 = csr_addr_i[1] | csr_addr_i[0];
  assign N388 = N1860 | N385;
  assign N389 = N386 | N387;
  assign N390 = N5410 | N388;
  assign N391 = N390 | N389;
  assign N393 = csr_addr_i[5] | csr_addr_i[4];
  assign N394 = csr_addr_i[3] | N280;
  assign N395 = csr_addr_i[1] | N170;
  assign N396 = N1860 | N393;
  assign N397 = N394 | N395;
  assign N398 = N5410 | N396;
  assign N399 = N398 | N397;
  assign N401 = csr_addr_i[5] | csr_addr_i[4];
  assign N402 = csr_addr_i[3] | N280;
  assign N403 = N180 | csr_addr_i[0];
  assign N404 = N1860 | N401;
  assign N405 = N402 | N403;
  assign N406 = N5410 | N404;
  assign N407 = N406 | N405;
  assign N409 = csr_addr_i[5] | csr_addr_i[4];
  assign N410 = csr_addr_i[3] | csr_addr_i[2];
  assign N411 = csr_addr_i[1] | csr_addr_i[0];
  assign N412 = N5419 | N409;
  assign N413 = N410 | N411;
  assign N414 = N5410 | N412;
  assign N415 = N414 | N413;
  assign N417 = csr_addr_i[5] | csr_addr_i[4];
  assign N418 = csr_addr_i[3] | csr_addr_i[2];
  assign N419 = csr_addr_i[1] | N170;
  assign N420 = N5419 | N417;
  assign N421 = N418 | N419;
  assign N422 = N5410 | N420;
  assign N423 = N422 | N421;
  assign N425 = csr_addr_i[5] | csr_addr_i[4];
  assign N426 = csr_addr_i[3] | csr_addr_i[2];
  assign N427 = N180 | csr_addr_i[0];
  assign N428 = N5419 | N425;
  assign N429 = N426 | N427;
  assign N430 = N5410 | N428;
  assign N431 = N430 | N429;
  assign N433 = csr_addr_i[5] | csr_addr_i[4];
  assign N434 = csr_addr_i[3] | csr_addr_i[2];
  assign N435 = N180 | N170;
  assign N436 = N5419 | N433;
  assign N437 = N434 | N435;
  assign N438 = N5410 | N436;
  assign N439 = N438 | N437;
  assign N441 = csr_addr_i[5] | csr_addr_i[4];
  assign N442 = csr_addr_i[3] | N280;
  assign N443 = csr_addr_i[1] | csr_addr_i[0];
  assign N444 = N5419 | N441;
  assign N445 = N442 | N443;
  assign N446 = N5410 | N444;
  assign N447 = N446 | N445;
  assign N449 = csr_addr_i[5] | N5553;
  assign N450 = csr_addr_i[3] | csr_addr_i[2];
  assign N451 = csr_addr_i[1] | N170;
  assign N452 = N1858 | N5406;
  assign N453 = N1860 | N449;
  assign N454 = N450 | N451;
  assign N455 = N452 | N453;
  assign N456 = N455 | N454;
  assign N458 = csr_addr_i[5] | N5553;
  assign N459 = csr_addr_i[3] | csr_addr_i[2];
  assign N460 = N180 | csr_addr_i[0];
  assign N461 = N1860 | N458;
  assign N462 = N459 | N460;
  assign N463 = N452 | N461;
  assign N464 = N463 | N462;
  assign N466 = csr_addr_i[5] | N5553;
  assign N467 = csr_addr_i[3] | csr_addr_i[2];
  assign N468 = N180 | N170;
  assign N469 = N1860 | N466;
  assign N470 = N467 | N468;
  assign N471 = N452 | N469;
  assign N472 = N471 | N470;
  assign N474 = csr_addr_i[5] | N5553;
  assign N475 = csr_addr_i[3] | N280;
  assign N476 = csr_addr_i[1] | csr_addr_i[0];
  assign N477 = N1860 | N474;
  assign N478 = N475 | N476;
  assign N479 = N452 | N477;
  assign N480 = N479 | N478;
  assign N482 = csr_addr_i[5] | csr_addr_i[4];
  assign N483 = csr_addr_i[3] | csr_addr_i[2];
  assign N484 = csr_addr_i[1] | csr_addr_i[0];
  assign N485 = N197 | N5406;
  assign N486 = N1860 | N482;
  assign N487 = N483 | N484;
  assign N488 = N485 | N486;
  assign N489 = N488 | N487;
  assign N491 = csr_addr_i[5] | csr_addr_i[4];
  assign N492 = csr_addr_i[3] | csr_addr_i[2];
  assign N493 = N180 | csr_addr_i[0];
  assign N494 = N1860 | N491;
  assign N495 = N492 | N493;
  assign N496 = N485 | N494;
  assign N497 = N496 | N495;
  assign N499 = csr_addr_i[5] | csr_addr_i[4];
  assign N500 = csr_addr_i[3] | csr_addr_i[2];
  assign N501 = csr_addr_i[1] | N170;
  assign N502 = N1860 | N499;
  assign N503 = N500 | N501;
  assign N504 = N1851 | N502;
  assign N505 = N504 | N503;
  assign N507 = csr_addr_i[5] | csr_addr_i[4];
  assign N508 = csr_addr_i[3] | csr_addr_i[2];
  assign N509 = csr_addr_i[1] | csr_addr_i[0];
  assign N510 = N1860 | N507;
  assign N511 = N508 | N509;
  assign N512 = N1851 | N510;
  assign N513 = N512 | N511;
  assign N515 = csr_addr_i[5] | csr_addr_i[4];
  assign N516 = csr_addr_i[3] | csr_addr_i[2];
  assign N517 = csr_addr_i[1] | csr_addr_i[0];
  assign N518 = N1860 | N515;
  assign N519 = N516 | N517;
  assign N520 = N1864 | N518;
  assign N521 = N520 | N519;
  assign N523 = csr_addr_i[5] | csr_addr_i[4];
  assign N524 = csr_addr_i[3] | csr_addr_i[2];
  assign N525 = N180 | csr_addr_i[0];
  assign N526 = N1860 | N523;
  assign N527 = N524 | N525;
  assign N528 = N1864 | N526;
  assign N529 = N528 | N527;
  assign N531 = csr_addr_i[5] | csr_addr_i[4];
  assign N532 = csr_addr_i[3] | csr_addr_i[2];
  assign N533 = N180 | N170;
  assign N534 = N1860 | N531;
  assign N535 = N532 | N533;
  assign N536 = N1864 | N534;
  assign N537 = N536 | N535;
  assign N538 = csr_addr_i[5] | csr_addr_i[4];
  assign N539 = csr_addr_i[3] | N280;
  assign N540 = csr_addr_i[1] | csr_addr_i[0];
  assign N541 = N1860 | N538;
  assign N542 = N539 | N540;
  assign N543 = N1864 | N541;
  assign N544 = N543 | N542;
  assign N545 = csr_addr_i[5] | csr_addr_i[4];
  assign N546 = csr_addr_i[3] | N280;
  assign N547 = csr_addr_i[1] | N170;
  assign N548 = N1860 | N545;
  assign N549 = N546 | N547;
  assign N550 = N1864 | N548;
  assign N551 = N550 | N549;
  assign N552 = csr_addr_i[5] | csr_addr_i[4];
  assign N553 = csr_addr_i[3] | N280;
  assign N554 = N180 | csr_addr_i[0];
  assign N555 = N1860 | N552;
  assign N556 = N553 | N554;
  assign N557 = N1864 | N555;
  assign N558 = N557 | N556;
  assign N559 = csr_addr_i[5] | csr_addr_i[4];
  assign N560 = csr_addr_i[3] | N280;
  assign N561 = N180 | N170;
  assign N562 = N1860 | N559;
  assign N563 = N560 | N561;
  assign N564 = N1864 | N562;
  assign N565 = N564 | N563;
  assign N567 = csr_addr_i[5] | csr_addr_i[4];
  assign N568 = N566 | csr_addr_i[2];
  assign N569 = csr_addr_i[1] | csr_addr_i[0];
  assign N570 = N1860 | N567;
  assign N571 = N568 | N569;
  assign N572 = N1864 | N570;
  assign N573 = N572 | N571;
  assign N574 = csr_addr_i[5] | csr_addr_i[4];
  assign N575 = N566 | csr_addr_i[2];
  assign N576 = csr_addr_i[1] | N170;
  assign N577 = N1860 | N574;
  assign N578 = N575 | N576;
  assign N579 = N1864 | N577;
  assign N580 = N579 | N578;
  assign N581 = csr_addr_i[5] | csr_addr_i[4];
  assign N582 = N566 | csr_addr_i[2];
  assign N583 = N180 | csr_addr_i[0];
  assign N584 = N1860 | N581;
  assign N585 = N582 | N583;
  assign N586 = N1864 | N584;
  assign N587 = N586 | N585;
  assign N588 = csr_addr_i[5] | csr_addr_i[4];
  assign N589 = N566 | csr_addr_i[2];
  assign N590 = N180 | N170;
  assign N591 = N1860 | N588;
  assign N592 = N589 | N590;
  assign N593 = N1864 | N591;
  assign N594 = N593 | N592;
  assign N595 = csr_addr_i[5] | csr_addr_i[4];
  assign N596 = N566 | N280;
  assign N597 = csr_addr_i[1] | csr_addr_i[0];
  assign N598 = N1860 | N595;
  assign N599 = N596 | N597;
  assign N600 = N1864 | N598;
  assign N601 = N600 | N599;
  assign N602 = csr_addr_i[5] | csr_addr_i[4];
  assign N603 = N566 | N280;
  assign N604 = csr_addr_i[1] | N170;
  assign N605 = N1860 | N602;
  assign N606 = N603 | N604;
  assign N607 = N1864 | N605;
  assign N608 = N607 | N606;
  assign N609 = csr_addr_i[5] | csr_addr_i[4];
  assign N610 = N566 | N280;
  assign N611 = N180 | csr_addr_i[0];
  assign N612 = N1860 | N609;
  assign N613 = N610 | N611;
  assign N614 = N1864 | N612;
  assign N615 = N614 | N613;
  assign N616 = csr_addr_i[5] | csr_addr_i[4];
  assign N617 = N566 | N280;
  assign N618 = N180 | N170;
  assign N619 = N1860 | N616;
  assign N620 = N617 | N618;
  assign N621 = N1864 | N619;
  assign N622 = N621 | N620;
  assign N623 = csr_addr_i[5] | N5553;
  assign N624 = csr_addr_i[3] | csr_addr_i[2];
  assign N625 = csr_addr_i[1] | csr_addr_i[0];
  assign N626 = N1860 | N623;
  assign N627 = N624 | N625;
  assign N628 = N1864 | N626;
  assign N629 = N628 | N627;
  assign N631 = csr_addr_i[9] & N5550;
  assign N632 = csr_addr_i[9] & csr_addr_i[3];
  assign N633 = csr_addr_i[10] & csr_addr_i[9];
  assign N634 = csr_addr_i[2] & csr_addr_i[0];
  assign N635 = N633 & N634;
  assign N636 = csr_addr_i[11] & csr_addr_i[5];
  assign N637 = N636 & csr_addr_i[0];
  assign N638 = N1857 & csr_addr_i[9];
  assign N639 = N5552 & csr_addr_i[4];
  assign N640 = N638 & N639;
  assign N641 = N640 & csr_addr_i[0];
  assign N642 = N5551 & csr_addr_i[5];
  assign N643 = N642 & csr_addr_i[0];
  assign N644 = csr_addr_i[7] & N5552;
  assign N645 = N644 & csr_addr_i[0];
  assign N646 = csr_addr_i[2] & csr_addr_i[1];
  assign N647 = N633 & N646;
  assign N648 = N636 & csr_addr_i[1];
  assign N649 = N642 & csr_addr_i[1];
  assign N650 = N1857 & csr_addr_i[10];
  assign N651 = N5552 & csr_addr_i[1];
  assign N652 = N650 & N651;
  assign N653 = N644 & csr_addr_i[1];
  assign N654 = N5551 & N5553;
  assign N655 = N633 & N654;
  assign N656 = N655 & csr_addr_i[1];
  assign N657 = N5552 & N5553;
  assign N658 = N633 & N657;
  assign N659 = N658 & csr_addr_i[1];
  assign N660 = N650 & csr_addr_i[2];
  assign N661 = csr_addr_i[5] & csr_addr_i[2];
  assign N662 = csr_addr_i[9] & N280;
  assign N663 = N180 & N170;
  assign N664 = N676 & N662;
  assign N665 = N664 & N663;
  assign N666 = csr_addr_i[9] & N5551;
  assign N667 = csr_addr_i[4] & N280;
  assign N668 = N180 & N170;
  assign N669 = N666 & N667;
  assign N670 = N669 & N668;
  assign N671 = csr_addr_i[9] & N5552;
  assign N672 = csr_addr_i[4] & N280;
  assign N673 = N180 & N170;
  assign N674 = N671 & N672;
  assign N675 = N674 & N673;
  assign N676 = csr_addr_i[11] & csr_addr_i[10];
  assign N677 = csr_addr_i[9] & N5553;
  assign N678 = N676 & N677;
  assign N679 = N5553 & csr_addr_i[2];
  assign N680 = N633 & N679;
  assign N681 = N642 & N5553;
  assign N682 = csr_addr_i[9] & csr_addr_i[7];
  assign N683 = N5552 & N5553;
  assign N684 = N682 & N683;
  assign N685 = N5548 & csr_addr_i[9];
  assign N686 = N685 & csr_addr_i[7];
  assign N687 = N5548 & csr_addr_i[5];
  assign N688 = csr_addr_i[9] & csr_addr_i[2];
  assign N689 = csr_addr_i[1] & csr_addr_i[0];
  assign N690 = N688 & N689;
  assign N691 = N5549 & csr_addr_i[5];
  assign N692 = N650 & N5549;
  assign N693 = csr_addr_i[10] & N5549;
  assign N694 = N693 & csr_addr_i[8];
  assign N695 = N693 & csr_addr_i[7];
  assign N696 = csr_addr_i[10] & csr_addr_i[6];
  assign N697 = N5549 & csr_addr_i[4];
  assign N698 = N697 & csr_addr_i[1];
  assign N699 = N5549 & csr_addr_i[4];
  assign N700 = N699 & csr_addr_i[2];
  assign N701 = csr_addr_i[4] & csr_addr_i[3];
  assign N702 = N566 & N280;
  assign N703 = N180 & csr_addr_i[0];
  assign N704 = N693 & N702;
  assign N705 = N704 & N703;
  assign N706 = N5548 & csr_addr_i[4];
  assign N707 = N5548 & csr_addr_i[3];
  assign N708 = csr_addr_i[11] & N5548;
  assign N709 = N708 & csr_addr_i[0];
  assign N710 = N5549 & csr_addr_i[7];
  assign N711 = N710 & csr_addr_i[0];
  assign N712 = N5548 & csr_addr_i[2];
  assign N713 = csr_addr_i[1] & csr_addr_i[0];
  assign N714 = N712 & N713;
  assign N715 = N5549 & csr_addr_i[8];
  assign N716 = N5416 & csr_addr_i[1];
  assign N717 = N715 & N716;
  assign N718 = N717 & csr_addr_i[0];
  assign N719 = csr_addr_i[6] & csr_addr_i[2];
  assign N720 = N719 & csr_addr_i[0];
  assign N721 = N5416 & N280;
  assign N722 = N715 & N721;
  assign N723 = N722 & csr_addr_i[0];
  assign N724 = N5549 & csr_addr_i[1];
  assign N725 = N708 & N724;
  assign N726 = N710 & csr_addr_i[1];
  assign N727 = csr_addr_i[6] & csr_addr_i[2];
  assign N728 = N727 & csr_addr_i[1];
  assign N729 = N5416 & N280;
  assign N730 = N715 & N729;
  assign N731 = N730 & csr_addr_i[1];
  assign N732 = N708 & csr_addr_i[2];
  assign N733 = N5548 & N5550;
  assign N734 = N733 & csr_addr_i[2];
  assign N735 = csr_addr_i[7] & csr_addr_i[2];
  assign N736 = csr_addr_i[11] & csr_addr_i[6];
  assign N737 = N5550 & csr_addr_i[6];
  assign N738 = N710 & csr_addr_i[6];
  assign N739 = csr_addr_i[11] & N5549;
  assign N740 = N739 & csr_addr_i[7];
  assign N741 = N5550 & csr_addr_i[7];
  assign N742 = N739 & csr_addr_i[8];
  assign N743 = N1857 & N5550;
  assign N744 = N180 & N170;
  assign N745 = N743 & N744;
  assign N1551 = csr_addr_i[5] | csr_addr_i[4];
  assign N1552 = csr_addr_i[3] | csr_addr_i[2];
  assign N1553 = csr_addr_i[1] | N170;
  assign N1554 = N1860 | N1551;
  assign N1555 = N1552 | N1553;
  assign N1556 = N174 | N1554;
  assign N1557 = N1556 | N1555;
  assign N1559 = csr_addr_i[5] | csr_addr_i[4];
  assign N1560 = csr_addr_i[3] | csr_addr_i[2];
  assign N1561 = N180 | csr_addr_i[0];
  assign N1562 = N1860 | N1559;
  assign N1563 = N1560 | N1561;
  assign N1564 = N174 | N1562;
  assign N1565 = N1564 | N1563;
  assign N1567 = csr_addr_i[5] | csr_addr_i[4];
  assign N1568 = csr_addr_i[3] | csr_addr_i[2];
  assign N1569 = N180 | N170;
  assign N1570 = N1860 | N1567;
  assign N1571 = N1568 | N1569;
  assign N1572 = N174 | N1570;
  assign N1573 = N1572 | N1571;
  assign N1575 = csr_addr_i[5] | csr_addr_i[4];
  assign N1576 = csr_addr_i[3] | csr_addr_i[2];
  assign N1577 = csr_addr_i[1] | csr_addr_i[0];
  assign N1578 = N1860 | N1575;
  assign N1579 = N1576 | N1577;
  assign N1580 = N201 | N1578;
  assign N1581 = N1580 | N1579;
  assign N1583 = N5552 | N5553;
  assign N1584 = csr_addr_i[3] | csr_addr_i[2];
  assign N1585 = csr_addr_i[1] | csr_addr_i[0];
  assign N1586 = N207 | N1583;
  assign N1587 = N1584 | N1585;
  assign N1588 = N1851 | N1586;
  assign N1589 = N1588 | N1587;
  assign N1591 = N5552 | N5553;
  assign N1592 = csr_addr_i[3] | csr_addr_i[2];
  assign N1593 = csr_addr_i[1] | N170;
  assign N1594 = N207 | N1591;
  assign N1595 = N1592 | N1593;
  assign N1596 = N1851 | N1594;
  assign N1597 = N1596 | N1595;
  assign N1599 = N5552 | N5553;
  assign N1600 = csr_addr_i[3] | csr_addr_i[2];
  assign N1601 = N180 | csr_addr_i[0];
  assign N1602 = N207 | N1599;
  assign N1603 = N1600 | N1601;
  assign N1604 = N1851 | N1602;
  assign N1605 = N1604 | N1603;
  assign N1607 = N5552 | N5553;
  assign N1608 = csr_addr_i[3] | csr_addr_i[2];
  assign N1609 = N180 | N170;
  assign N1610 = N207 | N1607;
  assign N1611 = N1608 | N1609;
  assign N1612 = N1851 | N1610;
  assign N1613 = N1612 | N1611;
  assign N1615 = N5552 | csr_addr_i[4];
  assign N1616 = csr_addr_i[3] | csr_addr_i[2];
  assign N1617 = csr_addr_i[1] | csr_addr_i[0];
  assign N1618 = N207 | N1615;
  assign N1619 = N1616 | N1617;
  assign N1620 = N1851 | N1618;
  assign N1621 = N1620 | N1619;
  assign N1623 = N5552 | csr_addr_i[4];
  assign N1624 = csr_addr_i[3] | csr_addr_i[2];
  assign N1625 = csr_addr_i[1] | N170;
  assign N1626 = N207 | N1623;
  assign N1627 = N1624 | N1625;
  assign N1628 = N1851 | N1626;
  assign N1629 = N1628 | N1627;
  assign N1631 = N5552 | csr_addr_i[4];
  assign N1632 = csr_addr_i[3] | csr_addr_i[2];
  assign N1633 = N180 | csr_addr_i[0];
  assign N1634 = N207 | N1631;
  assign N1635 = N1632 | N1633;
  assign N1636 = N1851 | N1634;
  assign N1637 = N1636 | N1635;
  assign N1639 = N5552 | csr_addr_i[4];
  assign N1640 = csr_addr_i[3] | csr_addr_i[2];
  assign N1641 = N180 | N170;
  assign N1642 = N207 | N1639;
  assign N1643 = N1640 | N1641;
  assign N1644 = N1851 | N1642;
  assign N1645 = N1644 | N1643;
  assign N1647 = csr_addr_i[5] | csr_addr_i[4];
  assign N1648 = csr_addr_i[3] | csr_addr_i[2];
  assign N1649 = csr_addr_i[1] | csr_addr_i[0];
  assign N1650 = N1860 | N1647;
  assign N1651 = N1648 | N1649;
  assign N1652 = N5423 | N1650;
  assign N1653 = N1652 | N1651;
  assign N1655 = csr_addr_i[5] | csr_addr_i[4];
  assign N1656 = csr_addr_i[3] | N280;
  assign N1657 = csr_addr_i[1] | csr_addr_i[0];
  assign N1658 = N1860 | N1655;
  assign N1659 = N1656 | N1657;
  assign N1660 = N5423 | N1658;
  assign N1661 = N1660 | N1659;
  assign N1663 = csr_addr_i[5] | csr_addr_i[4];
  assign N1664 = csr_addr_i[3] | N280;
  assign N1665 = csr_addr_i[1] | csr_addr_i[0];
  assign N1666 = N5419 | N1663;
  assign N1667 = N1664 | N1665;
  assign N1668 = N5423 | N1666;
  assign N1669 = N1668 | N1667;
  assign N1671 = csr_addr_i[5] | csr_addr_i[4];
  assign N1672 = csr_addr_i[3] | N280;
  assign N1673 = N180 | csr_addr_i[0];
  assign N1674 = N1860 | N1671;
  assign N1675 = N1672 | N1673;
  assign N1676 = N5423 | N1674;
  assign N1677 = N1676 | N1675;
  assign N1679 = csr_addr_i[5] | csr_addr_i[4];
  assign N1680 = csr_addr_i[3] | N280;
  assign N1681 = csr_addr_i[1] | N170;
  assign N1682 = N1860 | N1679;
  assign N1683 = N1680 | N1681;
  assign N1684 = N5423 | N1682;
  assign N1685 = N1684 | N1683;
  assign N1687 = csr_addr_i[5] | csr_addr_i[4];
  assign N1688 = csr_addr_i[3] | csr_addr_i[2];
  assign N1689 = csr_addr_i[1] | csr_addr_i[0];
  assign N1690 = N5419 | N1687;
  assign N1691 = N1688 | N1689;
  assign N1692 = N5423 | N1690;
  assign N1693 = N1692 | N1691;
  assign N1695 = csr_addr_i[5] | csr_addr_i[4];
  assign N1696 = csr_addr_i[3] | csr_addr_i[2];
  assign N1697 = csr_addr_i[1] | N170;
  assign N1698 = N5419 | N1695;
  assign N1699 = N1696 | N1697;
  assign N1700 = N5423 | N1698;
  assign N1701 = N1700 | N1699;
  assign N1703 = csr_addr_i[5] | csr_addr_i[4];
  assign N1704 = csr_addr_i[3] | csr_addr_i[2];
  assign N1705 = N180 | csr_addr_i[0];
  assign N1706 = N5419 | N1703;
  assign N1707 = N1704 | N1705;
  assign N1708 = N5423 | N1706;
  assign N1709 = N1708 | N1707;
  assign N1711 = csr_addr_i[5] | csr_addr_i[4];
  assign N1712 = csr_addr_i[3] | csr_addr_i[2];
  assign N1713 = N180 | N170;
  assign N1714 = N5419 | N1711;
  assign N1715 = N1712 | N1713;
  assign N1716 = N5423 | N1714;
  assign N1717 = N1716 | N1715;
  assign N1719 = csr_addr_i[5] | csr_addr_i[4];
  assign N1720 = csr_addr_i[3] | csr_addr_i[2];
  assign N1721 = csr_addr_i[1] | csr_addr_i[0];
  assign N1722 = N207 | N1719;
  assign N1723 = N1720 | N1721;
  assign N1724 = N5423 | N1722;
  assign N1725 = N1724 | N1723;
  assign N1727 = csr_addr_i[5] | csr_addr_i[4];
  assign N1728 = csr_addr_i[3] | csr_addr_i[2];
  assign N1729 = csr_addr_i[1] | csr_addr_i[0];
  assign N1730 = N1860 | N1727;
  assign N1731 = N1728 | N1729;
  assign N1732 = N5410 | N1730;
  assign N1733 = N1732 | N1731;
  assign N1735 = csr_addr_i[5] | csr_addr_i[4];
  assign N1736 = csr_addr_i[3] | csr_addr_i[2];
  assign N1737 = csr_addr_i[1] | N170;
  assign N1738 = N1860 | N1735;
  assign N1739 = N1736 | N1737;
  assign N1740 = N5410 | N1738;
  assign N1741 = N1740 | N1739;
  assign N1743 = csr_addr_i[5] | csr_addr_i[4];
  assign N1744 = csr_addr_i[3] | csr_addr_i[2];
  assign N1745 = N180 | csr_addr_i[0];
  assign N1746 = N1860 | N1743;
  assign N1747 = N1744 | N1745;
  assign N1748 = N5410 | N1746;
  assign N1749 = N1748 | N1747;
  assign N1751 = csr_addr_i[5] | csr_addr_i[4];
  assign N1752 = csr_addr_i[3] | csr_addr_i[2];
  assign N1753 = N180 | N170;
  assign N1754 = N1860 | N1751;
  assign N1755 = N1752 | N1753;
  assign N1756 = N5410 | N1754;
  assign N1757 = N1756 | N1755;
  assign N1759 = csr_addr_i[5] | csr_addr_i[4];
  assign N1760 = csr_addr_i[3] | N280;
  assign N1761 = csr_addr_i[1] | csr_addr_i[0];
  assign N1762 = N1860 | N1759;
  assign N1763 = N1760 | N1761;
  assign N1764 = N5410 | N1762;
  assign N1765 = N1764 | N1763;
  assign N1767 = csr_addr_i[5] | csr_addr_i[4];
  assign N1768 = csr_addr_i[3] | N280;
  assign N1769 = csr_addr_i[1] | N170;
  assign N1770 = N1860 | N1767;
  assign N1771 = N1768 | N1769;
  assign N1772 = N5410 | N1770;
  assign N1773 = N1772 | N1771;
  assign N1775 = csr_addr_i[5] | csr_addr_i[4];
  assign N1776 = csr_addr_i[3] | N280;
  assign N1777 = N180 | csr_addr_i[0];
  assign N1778 = N1860 | N1775;
  assign N1779 = N1776 | N1777;
  assign N1780 = N5410 | N1778;
  assign N1781 = N1780 | N1779;
  assign N1783 = csr_addr_i[5] | csr_addr_i[4];
  assign N1784 = csr_addr_i[3] | csr_addr_i[2];
  assign N1785 = csr_addr_i[1] | csr_addr_i[0];
  assign N1786 = N5419 | N1783;
  assign N1787 = N1784 | N1785;
  assign N1788 = N5410 | N1786;
  assign N1789 = N1788 | N1787;
  assign N1791 = csr_addr_i[5] | csr_addr_i[4];
  assign N1792 = csr_addr_i[3] | csr_addr_i[2];
  assign N1793 = csr_addr_i[1] | N170;
  assign N1794 = N5419 | N1791;
  assign N1795 = N1792 | N1793;
  assign N1796 = N5410 | N1794;
  assign N1797 = N1796 | N1795;
  assign N1799 = csr_addr_i[5] | csr_addr_i[4];
  assign N1800 = csr_addr_i[3] | csr_addr_i[2];
  assign N1801 = N180 | csr_addr_i[0];
  assign N1802 = N5419 | N1799;
  assign N1803 = N1800 | N1801;
  assign N1804 = N5410 | N1802;
  assign N1805 = N1804 | N1803;
  assign N1807 = csr_addr_i[5] | csr_addr_i[4];
  assign N1808 = csr_addr_i[3] | csr_addr_i[2];
  assign N1809 = N180 | N170;
  assign N1810 = N5419 | N1807;
  assign N1811 = N1808 | N1809;
  assign N1812 = N5410 | N1810;
  assign N1813 = N1812 | N1811;
  assign N1815 = csr_addr_i[5] | csr_addr_i[4];
  assign N1816 = csr_addr_i[3] | N280;
  assign N1817 = csr_addr_i[1] | csr_addr_i[0];
  assign N1818 = N5419 | N1815;
  assign N1819 = N1816 | N1817;
  assign N1820 = N5410 | N1818;
  assign N1821 = N1820 | N1819;
  assign N1823 = csr_addr_i[5] | csr_addr_i[4];
  assign N1824 = csr_addr_i[3] | csr_addr_i[2];
  assign N1825 = csr_addr_i[1] | csr_addr_i[0];
  assign N1826 = N1860 | N1823;
  assign N1827 = N1824 | N1825;
  assign N1828 = N485 | N1826;
  assign N1829 = N1828 | N1827;
  assign N1831 = csr_addr_i[5] | csr_addr_i[4];
  assign N1832 = csr_addr_i[3] | csr_addr_i[2];
  assign N1833 = N180 | csr_addr_i[0];
  assign N1834 = N1860 | N1831;
  assign N1835 = N1832 | N1833;
  assign N1836 = N485 | N1834;
  assign N1837 = N1836 | N1835;
  assign N1839 = csr_addr_i[5] | csr_addr_i[4];
  assign N1840 = csr_addr_i[3] | csr_addr_i[2];
  assign N1841 = csr_addr_i[1] | N170;
  assign N1842 = N1860 | N1839;
  assign N1843 = N1840 | N1841;
  assign N1844 = N1851 | N1842;
  assign N1845 = N1844 | N1843;
  assign N1847 = csr_addr_i[11] | N5548;
  assign N1848 = csr_addr_i[5] | csr_addr_i[4];
  assign N1849 = csr_addr_i[3] | csr_addr_i[2];
  assign N1850 = csr_addr_i[1] | csr_addr_i[0];
  assign N1851 = N1847 | N5406;
  assign N1852 = N1860 | N1848;
  assign N1853 = N1849 | N1850;
  assign N1854 = N1851 | N1852;
  assign N1855 = N1854 | N1853;
  assign N1858 = N1857 | N5548;
  assign N1859 = csr_addr_i[9] | csr_addr_i[8];
  assign N1860 = csr_addr_i[7] | csr_addr_i[6];
  assign N1861 = csr_addr_i[5] | csr_addr_i[4];
  assign N1862 = csr_addr_i[3] | csr_addr_i[2];
  assign N1863 = N180 | N170;
  assign N1864 = N1858 | N1859;
  assign N1865 = N1860 | N1861;
  assign N1866 = N1862 | N1863;
  assign N1867 = N1864 | N1865;
  assign N1868 = N1867 | N1866;
  assign N1869 = csr_addr_i[5] | csr_addr_i[4];
  assign N1870 = csr_addr_i[3] | N280;
  assign N1871 = csr_addr_i[1] | csr_addr_i[0];
  assign N1872 = N1860 | N1869;
  assign N1873 = N1870 | N1871;
  assign N1874 = N1864 | N1872;
  assign N1875 = N1874 | N1873;
  assign N1876 = csr_addr_i[5] | csr_addr_i[4];
  assign N1877 = csr_addr_i[3] | N280;
  assign N1878 = csr_addr_i[1] | N170;
  assign N1879 = N1860 | N1876;
  assign N1880 = N1877 | N1878;
  assign N1881 = N1864 | N1879;
  assign N1882 = N1881 | N1880;
  assign N1883 = csr_addr_i[5] | csr_addr_i[4];
  assign N1884 = csr_addr_i[3] | N280;
  assign N1885 = N180 | csr_addr_i[0];
  assign N1886 = N1860 | N1883;
  assign N1887 = N1884 | N1885;
  assign N1888 = N1864 | N1886;
  assign N1889 = N1888 | N1887;
  assign N1890 = csr_addr_i[5] | csr_addr_i[4];
  assign N1891 = csr_addr_i[3] | N280;
  assign N1892 = N180 | N170;
  assign N1893 = N1860 | N1890;
  assign N1894 = N1891 | N1892;
  assign N1895 = N1864 | N1893;
  assign N1896 = N1895 | N1894;
  assign N1897 = csr_addr_i[5] | csr_addr_i[4];
  assign N1898 = N566 | csr_addr_i[2];
  assign N1899 = csr_addr_i[1] | csr_addr_i[0];
  assign N1900 = N1860 | N1897;
  assign N1901 = N1898 | N1899;
  assign N1902 = N1864 | N1900;
  assign N1903 = N1902 | N1901;
  assign N1904 = csr_addr_i[5] | csr_addr_i[4];
  assign N1905 = N566 | csr_addr_i[2];
  assign N1906 = csr_addr_i[1] | N170;
  assign N1907 = N1860 | N1904;
  assign N1908 = N1905 | N1906;
  assign N1909 = N1864 | N1907;
  assign N1910 = N1909 | N1908;
  assign N1911 = csr_addr_i[5] | csr_addr_i[4];
  assign N1912 = N566 | csr_addr_i[2];
  assign N1913 = N180 | csr_addr_i[0];
  assign N1914 = N1860 | N1911;
  assign N1915 = N1912 | N1913;
  assign N1916 = N1864 | N1914;
  assign N1917 = N1916 | N1915;
  assign N1918 = csr_addr_i[5] | csr_addr_i[4];
  assign N1919 = N566 | csr_addr_i[2];
  assign N1920 = N180 | N170;
  assign N1921 = N1860 | N1918;
  assign N1922 = N1919 | N1920;
  assign N1923 = N1864 | N1921;
  assign N1924 = N1923 | N1922;
  assign N1925 = csr_addr_i[5] | csr_addr_i[4];
  assign N1926 = N566 | N280;
  assign N1927 = csr_addr_i[1] | csr_addr_i[0];
  assign N1928 = N1860 | N1925;
  assign N1929 = N1926 | N1927;
  assign N1930 = N1864 | N1928;
  assign N1931 = N1930 | N1929;
  assign N1932 = csr_addr_i[5] | csr_addr_i[4];
  assign N1933 = N566 | N280;
  assign N1934 = csr_addr_i[1] | N170;
  assign N1935 = N1860 | N1932;
  assign N1936 = N1933 | N1934;
  assign N1937 = N1864 | N1935;
  assign N1938 = N1937 | N1936;
  assign N1939 = csr_addr_i[5] | csr_addr_i[4];
  assign N1940 = N566 | N280;
  assign N1941 = N180 | csr_addr_i[0];
  assign N1942 = N1860 | N1939;
  assign N1943 = N1940 | N1941;
  assign N1944 = N1864 | N1942;
  assign N1945 = N1944 | N1943;
  assign N4156 = (N4092)? mideleg_d[0] : 
                 (N4094)? mideleg_q_1 : 
                 (N4096)? mideleg_d[2] : 
                 (N4098)? mideleg_d[3] : 
                 (N4100)? mideleg_d[4] : 
                 (N4102)? mideleg_q_5 : 
                 (N4104)? mideleg_d[6] : 
                 (N4106)? mideleg_d[7] : 
                 (N4108)? mideleg_d[8] : 
                 (N4110)? mideleg_q[9] : 
                 (N4112)? mideleg_d[10] : 
                 (N4114)? mideleg_d[11] : 
                 (N4116)? mideleg_d[12] : 
                 (N4118)? mideleg_d[13] : 
                 (N4120)? mideleg_d[14] : 
                 (N4122)? mideleg_d[15] : 
                 (N4124)? mideleg_d[16] : 
                 (N4126)? mideleg_d[17] : 
                 (N4128)? mideleg_d[18] : 
                 (N4130)? mideleg_d[19] : 
                 (N4132)? mideleg_d[20] : 
                 (N4134)? mideleg_d[21] : 
                 (N4136)? mideleg_d[22] : 
                 (N4138)? mideleg_d[23] : 
                 (N4140)? mideleg_d[24] : 
                 (N4142)? mideleg_d[25] : 
                 (N4144)? mideleg_d[26] : 
                 (N4146)? mideleg_d[27] : 
                 (N4148)? mideleg_d[28] : 
                 (N4150)? mideleg_d[29] : 
                 (N4152)? mideleg_d[30] : 
                 (N4154)? mideleg_d[31] : 
                 (N4093)? mideleg_d[32] : 
                 (N4095)? mideleg_d[33] : 
                 (N4097)? mideleg_d[34] : 
                 (N4099)? mideleg_d[35] : 
                 (N4101)? mideleg_d[36] : 
                 (N4103)? mideleg_d[37] : 
                 (N4105)? mideleg_d[38] : 
                 (N4107)? mideleg_d[39] : 
                 (N4109)? mideleg_d[40] : 
                 (N4111)? mideleg_d[41] : 
                 (N4113)? mideleg_d[42] : 
                 (N4115)? mideleg_d[43] : 
                 (N4117)? mideleg_d[44] : 
                 (N4119)? mideleg_d[45] : 
                 (N4121)? mideleg_d[46] : 
                 (N4123)? mideleg_d[47] : 
                 (N4125)? mideleg_d[48] : 
                 (N4127)? mideleg_d[49] : 
                 (N4129)? mideleg_d[50] : 
                 (N4131)? mideleg_d[51] : 
                 (N4133)? mideleg_d[52] : 
                 (N4135)? mideleg_d[53] : 
                 (N4137)? mideleg_d[54] : 
                 (N4139)? mideleg_d[55] : 
                 (N4141)? mideleg_d[56] : 
                 (N4143)? mideleg_d[57] : 
                 (N4145)? mideleg_d[58] : 
                 (N4147)? mideleg_d[59] : 
                 (N4149)? mideleg_d[60] : 
                 (N4151)? mideleg_d[61] : 
                 (N4153)? mideleg_d[62] : 
                 (N4155)? mideleg_d[63] : 1'b0;
  assign N4157 = (N4092)? medeleg_q_0 : 
                 (N4094)? medeleg_d[1] : 
                 (N4096)? medeleg_d[2] : 
                 (N4098)? medeleg_q_3 : 
                 (N4100)? medeleg_d[4] : 
                 (N4102)? medeleg_d[5] : 
                 (N4104)? medeleg_d[6] : 
                 (N4106)? medeleg_d[7] : 
                 (N4108)? medeleg_q_8 : 
                 (N4110)? medeleg_d[9] : 
                 (N4112)? medeleg_d[10] : 
                 (N4114)? medeleg_d[11] : 
                 (N4116)? medeleg_q[12] : 
                 (N4118)? medeleg_q[13] : 
                 (N4120)? medeleg_d[14] : 
                 (N4122)? medeleg_q_15 : 
                 (N4124)? medeleg_d[16] : 
                 (N4126)? medeleg_d[17] : 
                 (N4128)? medeleg_d[18] : 
                 (N4130)? medeleg_d[19] : 
                 (N4132)? medeleg_d[20] : 
                 (N4134)? medeleg_d[21] : 
                 (N4136)? medeleg_d[22] : 
                 (N4138)? medeleg_d[23] : 
                 (N4140)? medeleg_d[24] : 
                 (N4142)? medeleg_d[25] : 
                 (N4144)? medeleg_d[26] : 
                 (N4146)? medeleg_d[27] : 
                 (N4148)? medeleg_d[28] : 
                 (N4150)? medeleg_d[29] : 
                 (N4152)? medeleg_d[30] : 
                 (N4154)? medeleg_d[31] : 
                 (N4093)? medeleg_d[32] : 
                 (N4095)? medeleg_d[33] : 
                 (N4097)? medeleg_d[34] : 
                 (N4099)? medeleg_d[35] : 
                 (N4101)? medeleg_d[36] : 
                 (N4103)? medeleg_d[37] : 
                 (N4105)? medeleg_d[38] : 
                 (N4107)? medeleg_d[39] : 
                 (N4109)? medeleg_d[40] : 
                 (N4111)? medeleg_d[41] : 
                 (N4113)? medeleg_d[42] : 
                 (N4115)? medeleg_d[43] : 
                 (N4117)? medeleg_d[44] : 
                 (N4119)? medeleg_d[45] : 
                 (N4121)? medeleg_d[46] : 
                 (N4123)? medeleg_d[47] : 
                 (N4125)? medeleg_d[48] : 
                 (N4127)? medeleg_d[49] : 
                 (N4129)? medeleg_d[50] : 
                 (N4131)? medeleg_d[51] : 
                 (N4133)? medeleg_d[52] : 
                 (N4135)? medeleg_d[53] : 
                 (N4137)? medeleg_d[54] : 
                 (N4139)? medeleg_d[55] : 
                 (N4141)? medeleg_d[56] : 
                 (N4143)? medeleg_d[57] : 
                 (N4145)? medeleg_d[58] : 
                 (N4147)? medeleg_d[59] : 
                 (N4149)? medeleg_d[60] : 
                 (N4151)? medeleg_d[61] : 
                 (N4153)? medeleg_d[62] : 
                 (N4155)? medeleg_d[63] : 1'b0;
  assign N4564 = priv_lvl_o[1] & priv_lvl_o[0];
  assign N4565 = priv_lvl_o[1] | N5543;
  assign N4568 = N4567 & N5543;
  assign N4569 = N4567 | priv_lvl_o[0];
  assign N4933 = N4945 | N4954;
  assign N4935 = N4941 | N4960;
  assign N4938 = N4937 | csr_op_i[4];
  assign N4939 = csr_op_i[3] | csr_op_i[2];
  assign N4940 = csr_op_i[1] | N4948;
  assign N4941 = N4938 | N4939;
  assign N4942 = N4941 | N4940;
  assign N4944 = N5512 | N4952;
  assign N4945 = N4958 | N4944;
  assign N4946 = N4945 | N4949;
  assign N4949 = N5513 | N4948;
  assign N4950 = N4955 | N4949;
  assign N4953 = csr_op_i[3] | N4952;
  assign N4954 = N5513 | csr_op_i[0];
  assign N4955 = N4958 | N4953;
  assign N4956 = N4955 | N4954;
  assign N4958 = csr_op_i[5] | N5511;
  assign N4959 = N5512 | csr_op_i[2];
  assign N4960 = csr_op_i[1] | csr_op_i[0];
  assign N4961 = N4958 | N4959;
  assign N4962 = N4961 | N4960;
  assign N5233 = (N5217)? mideleg_d[0] : 
                 (N5219)? mideleg_q_1 : 
                 (N5221)? mideleg_d[2] : 
                 (N5223)? mideleg_d[3] : 
                 (N5225)? mideleg_d[4] : 
                 (N5227)? mideleg_q_5 : 
                 (N5229)? mideleg_d[6] : 
                 (N5231)? mideleg_d[7] : 
                 (N5218)? mideleg_d[8] : 
                 (N5220)? mideleg_q[9] : 
                 (N5222)? mideleg_d[10] : 
                 (N5224)? mideleg_d[11] : 
                 (N5226)? mideleg_d[12] : 
                 (N5228)? mideleg_d[13] : 
                 (N5230)? mideleg_d[14] : 
                 (N5232)? mideleg_d[15] : 
                 (N0)? mideleg_d[16] : 
                 (N0)? mideleg_d[17] : 
                 (N0)? mideleg_d[18] : 
                 (N0)? mideleg_d[19] : 
                 (N0)? mideleg_d[20] : 
                 (N0)? mideleg_d[21] : 
                 (N0)? mideleg_d[22] : 
                 (N0)? mideleg_d[23] : 
                 (N0)? mideleg_d[24] : 
                 (N0)? mideleg_d[25] : 
                 (N0)? mideleg_d[26] : 
                 (N0)? mideleg_d[27] : 
                 (N0)? mideleg_d[28] : 
                 (N0)? mideleg_d[29] : 
                 (N0)? mideleg_d[30] : 
                 (N0)? mideleg_d[31] : 
                 (N0)? mideleg_d[32] : 
                 (N0)? mideleg_d[33] : 
                 (N0)? mideleg_d[34] : 
                 (N0)? mideleg_d[35] : 
                 (N0)? mideleg_d[36] : 
                 (N0)? mideleg_d[37] : 
                 (N0)? mideleg_d[38] : 
                 (N0)? mideleg_d[39] : 
                 (N0)? mideleg_d[40] : 
                 (N0)? mideleg_d[41] : 
                 (N0)? mideleg_d[42] : 
                 (N0)? mideleg_d[43] : 
                 (N0)? mideleg_d[44] : 
                 (N0)? mideleg_d[45] : 
                 (N0)? mideleg_d[46] : 
                 (N0)? mideleg_d[47] : 
                 (N0)? mideleg_d[48] : 
                 (N0)? mideleg_d[49] : 
                 (N0)? mideleg_d[50] : 
                 (N0)? mideleg_d[51] : 
                 (N0)? mideleg_d[52] : 
                 (N0)? mideleg_d[53] : 
                 (N0)? mideleg_d[54] : 
                 (N0)? mideleg_d[55] : 
                 (N0)? mideleg_d[56] : 
                 (N0)? mideleg_d[57] : 
                 (N0)? mideleg_d[58] : 
                 (N0)? mideleg_d[59] : 
                 (N0)? mideleg_d[60] : 
                 (N0)? mideleg_d[61] : 
                 (N0)? mideleg_d[62] : 
                 (N0)? mideleg_d[63] : 1'b0;
  assign N0 = 1'b0;
  assign N5246 = { N5244, N5245 } != csr_addr_i[9:8];
  assign N5406 = N5549 | N5550;
  assign N5407 = csr_addr_i[5] | csr_addr_i[4];
  assign N5408 = csr_addr_i[3] | N280;
  assign N5409 = csr_addr_i[1] | csr_addr_i[0];
  assign N5410 = N5417 | N5406;
  assign N5411 = N5419 | N5407;
  assign N5412 = N5408 | N5409;
  assign N5413 = N5410 | N5411;
  assign N5414 = N5413 | N5412;
  assign N5417 = csr_addr_i[11] | csr_addr_i[10];
  assign N5418 = csr_addr_i[9] | N5550;
  assign N5419 = csr_addr_i[7] | N5416;
  assign N5420 = csr_addr_i[5] | csr_addr_i[4];
  assign N5421 = csr_addr_i[3] | N280;
  assign N5422 = csr_addr_i[1] | csr_addr_i[0];
  assign N5423 = N5417 | N5418;
  assign N5424 = N5419 | N5420;
  assign N5425 = N5421 | N5422;
  assign N5426 = N5423 | N5424;
  assign N5427 = N5426 | N5425;

  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      halt_csr_o <= 1'b0;
    end else if(N5269) begin
      halt_csr_o <= wfi_d;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      priv_lvl_q[1] <= 1'b1;
    end else if(1'b1) begin
      priv_lvl_q[1] <= priv_lvl_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      priv_lvl_q[0] <= 1'b1;
    end else if(1'b1) begin
      priv_lvl_q[0] <= priv_lvl_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[6] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[6] <= fcsr_d_fprec__6_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[5] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[5] <= fcsr_d_fprec__5_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[4] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[4] <= fcsr_d_fprec__4_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[3] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[3] <= fcsr_d_fprec__3_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[2] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[2] <= fcsr_d_fprec__2_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[1] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[1] <= fcsr_d_fprec__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fprec_o[0] <= 1'b0;
    end else if(1'b1) begin
      fprec_o[0] <= fcsr_d_fprec__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      frm_o[2] <= 1'b0;
    end else if(1'b1) begin
      frm_o[2] <= fcsr_d_frm__2_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      frm_o[1] <= 1'b0;
    end else if(1'b1) begin
      frm_o[1] <= fcsr_d_frm__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      frm_o[0] <= 1'b0;
    end else if(1'b1) begin
      frm_o[0] <= fcsr_d_frm__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fflags_o[4] <= 1'b0;
    end else if(1'b1) begin
      fflags_o[4] <= fcsr_d_fflags__4_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fflags_o[3] <= 1'b0;
    end else if(1'b1) begin
      fflags_o[3] <= fcsr_d_fflags__3_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fflags_o[2] <= 1'b0;
    end else if(1'b1) begin
      fflags_o[2] <= fcsr_d_fflags__2_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fflags_o[1] <= 1'b0;
    end else if(1'b1) begin
      fflags_o[1] <= fcsr_d_fflags__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fflags_o[0] <= 1'b0;
    end else if(1'b1) begin
      fflags_o[0] <= fcsr_d_fflags__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      debug_mode_o <= 1'b0;
    end else if(1'b1) begin
      debug_mode_o <= debug_mode_d;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_xdebugver__31_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__31_ <= dcsr_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_xdebugver__30_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__30_ <= dcsr_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_xdebugver__29_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__29_ <= dcsr_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_xdebugver__28_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__28_ <= dcsr_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__27_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__27_ <= dcsr_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__26_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__26_ <= dcsr_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__25_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__25_ <= dcsr_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__24_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__24_ <= dcsr_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__23_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__23_ <= dcsr_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__22_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__22_ <= dcsr_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__21_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__21_ <= dcsr_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__20_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__20_ <= dcsr_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__19_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__19_ <= dcsr_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__18_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__18_ <= dcsr_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__17_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__17_ <= dcsr_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero2__16_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__16_ <= dcsr_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_ebreakm_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_ebreakm_ <= dcsr_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero1_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero1_ <= dcsr_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_ebreaks_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_ebreaks_ <= dcsr_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_ebreaku_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_ebreaku_ <= dcsr_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_stepie_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stepie_ <= dcsr_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_stopcount_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stopcount_ <= dcsr_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_stoptime_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stoptime_ <= dcsr_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_cause__8_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__8_ <= dcsr_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_cause__7_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__7_ <= dcsr_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_cause__6_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__6_ <= dcsr_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_zero0_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero0_ <= dcsr_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_mprven_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_mprven_ <= dcsr_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_nmip_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_nmip_ <= dcsr_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      single_step_o <= 1'b0;
    end else if(1'b1) begin
      single_step_o <= dcsr_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_prv__1_ <= 1'b1;
    end else if(1'b1) begin
      dcsr_q_prv__1_ <= dcsr_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcsr_q_prv__0_ <= 1'b1;
    end else if(1'b1) begin
      dcsr_q_prv__0_ <= dcsr_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[63] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[63] <= dpc_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[62] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[62] <= dpc_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[61] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[61] <= dpc_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[60] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[60] <= dpc_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[59] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[59] <= dpc_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[58] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[58] <= dpc_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[57] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[57] <= dpc_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[56] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[56] <= dpc_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[55] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[55] <= dpc_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[54] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[54] <= dpc_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[53] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[53] <= dpc_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[52] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[52] <= dpc_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[51] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[51] <= dpc_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[50] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[50] <= dpc_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[49] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[49] <= dpc_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[48] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[48] <= dpc_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[47] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[47] <= dpc_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[46] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[46] <= dpc_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[45] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[45] <= dpc_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[44] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[44] <= dpc_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[43] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[43] <= dpc_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[42] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[42] <= dpc_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[41] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[41] <= dpc_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[40] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[40] <= dpc_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[39] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[39] <= dpc_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[38] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[38] <= dpc_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[37] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[37] <= dpc_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[36] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[36] <= dpc_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[35] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[35] <= dpc_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[34] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[34] <= dpc_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[33] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[33] <= dpc_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[32] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[32] <= dpc_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[31] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[31] <= dpc_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[30] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[30] <= dpc_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[29] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[29] <= dpc_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[28] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[28] <= dpc_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[27] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[27] <= dpc_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[26] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[26] <= dpc_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[25] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[25] <= dpc_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[24] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[24] <= dpc_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[23] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[23] <= dpc_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[22] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[22] <= dpc_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[21] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[21] <= dpc_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[20] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[20] <= dpc_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[19] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[19] <= dpc_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[18] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[18] <= dpc_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[17] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[17] <= dpc_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[16] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[16] <= dpc_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[15] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[15] <= dpc_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[14] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[14] <= dpc_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[13] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[13] <= dpc_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[12] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[12] <= dpc_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[11] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[11] <= dpc_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[10] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[10] <= dpc_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[9] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[9] <= dpc_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[8] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[8] <= dpc_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[7] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[7] <= dpc_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[6] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[6] <= dpc_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[5] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[5] <= dpc_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[4] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[4] <= dpc_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[3] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[3] <= dpc_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[2] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[2] <= dpc_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[1] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[1] <= dpc_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dpc_q[0] <= 1'b0;
    end else if(1'b1) begin
      dpc_q[0] <= dpc_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[63] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[63] <= dscratch0_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[62] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[62] <= dscratch0_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[61] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[61] <= dscratch0_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[60] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[60] <= dscratch0_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[59] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[59] <= dscratch0_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[58] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[58] <= dscratch0_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[57] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[57] <= dscratch0_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[56] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[56] <= dscratch0_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[55] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[55] <= dscratch0_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[54] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[54] <= dscratch0_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[53] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[53] <= dscratch0_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[52] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[52] <= dscratch0_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[51] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[51] <= dscratch0_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[50] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[50] <= dscratch0_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[49] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[49] <= dscratch0_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[48] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[48] <= dscratch0_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[47] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[47] <= dscratch0_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[46] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[46] <= dscratch0_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[45] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[45] <= dscratch0_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[44] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[44] <= dscratch0_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[43] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[43] <= dscratch0_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[42] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[42] <= dscratch0_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[41] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[41] <= dscratch0_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[40] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[40] <= dscratch0_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[39] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[39] <= dscratch0_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[38] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[38] <= dscratch0_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[37] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[37] <= dscratch0_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[36] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[36] <= dscratch0_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[35] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[35] <= dscratch0_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[34] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[34] <= dscratch0_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[33] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[33] <= dscratch0_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[32] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[32] <= dscratch0_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[31] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[31] <= dscratch0_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[30] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[30] <= dscratch0_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[29] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[29] <= dscratch0_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[28] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[28] <= dscratch0_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[27] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[27] <= dscratch0_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[26] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[26] <= dscratch0_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[25] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[25] <= dscratch0_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[24] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[24] <= dscratch0_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[23] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[23] <= dscratch0_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[22] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[22] <= dscratch0_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[21] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[21] <= dscratch0_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[20] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[20] <= dscratch0_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[19] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[19] <= dscratch0_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[18] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[18] <= dscratch0_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[17] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[17] <= dscratch0_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[16] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[16] <= dscratch0_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[15] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[15] <= dscratch0_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[14] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[14] <= dscratch0_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[13] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[13] <= dscratch0_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[12] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[12] <= dscratch0_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[11] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[11] <= dscratch0_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[10] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[10] <= dscratch0_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[9] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[9] <= dscratch0_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[8] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[8] <= dscratch0_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[7] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[7] <= dscratch0_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[6] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[6] <= dscratch0_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[5] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[5] <= dscratch0_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[4] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[4] <= dscratch0_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[3] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[3] <= dscratch0_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[2] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[2] <= dscratch0_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[1] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[1] <= dscratch0_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch0_q[0] <= 1'b0;
    end else if(1'b1) begin
      dscratch0_q[0] <= dscratch0_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[63] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[63] <= dscratch1_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[62] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[62] <= dscratch1_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[61] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[61] <= dscratch1_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[60] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[60] <= dscratch1_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[59] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[59] <= dscratch1_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[58] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[58] <= dscratch1_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[57] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[57] <= dscratch1_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[56] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[56] <= dscratch1_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[55] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[55] <= dscratch1_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[54] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[54] <= dscratch1_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[53] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[53] <= dscratch1_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[52] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[52] <= dscratch1_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[51] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[51] <= dscratch1_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[50] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[50] <= dscratch1_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[49] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[49] <= dscratch1_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[48] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[48] <= dscratch1_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[47] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[47] <= dscratch1_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[46] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[46] <= dscratch1_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[45] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[45] <= dscratch1_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[44] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[44] <= dscratch1_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[43] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[43] <= dscratch1_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[42] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[42] <= dscratch1_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[41] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[41] <= dscratch1_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[40] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[40] <= dscratch1_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[39] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[39] <= dscratch1_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[38] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[38] <= dscratch1_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[37] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[37] <= dscratch1_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[36] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[36] <= dscratch1_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[35] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[35] <= dscratch1_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[34] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[34] <= dscratch1_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[33] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[33] <= dscratch1_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[32] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[32] <= dscratch1_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[31] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[31] <= dscratch1_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[30] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[30] <= dscratch1_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[29] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[29] <= dscratch1_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[28] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[28] <= dscratch1_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[27] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[27] <= dscratch1_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[26] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[26] <= dscratch1_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[25] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[25] <= dscratch1_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[24] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[24] <= dscratch1_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[23] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[23] <= dscratch1_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[22] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[22] <= dscratch1_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[21] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[21] <= dscratch1_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[20] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[20] <= dscratch1_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[19] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[19] <= dscratch1_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[18] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[18] <= dscratch1_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[17] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[17] <= dscratch1_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[16] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[16] <= dscratch1_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[15] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[15] <= dscratch1_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[14] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[14] <= dscratch1_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[13] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[13] <= dscratch1_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[12] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[12] <= dscratch1_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[11] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[11] <= dscratch1_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[10] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[10] <= dscratch1_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[9] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[9] <= dscratch1_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[8] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[8] <= dscratch1_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[7] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[7] <= dscratch1_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[6] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[6] <= dscratch1_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[5] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[5] <= dscratch1_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[4] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[4] <= dscratch1_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[3] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[3] <= dscratch1_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[2] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[2] <= dscratch1_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[1] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[1] <= dscratch1_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dscratch1_q[0] <= 1'b0;
    end else if(1'b1) begin
      dscratch1_q[0] <= dscratch1_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_sd_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_sd_ <= mstatus_d_sd_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__62_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__62_ <= mstatus_d_wpri4__62_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__61_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__61_ <= mstatus_d_wpri4__61_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__60_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__60_ <= mstatus_d_wpri4__60_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__59_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__59_ <= mstatus_d_wpri4__59_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__58_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__58_ <= mstatus_d_wpri4__58_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__57_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__57_ <= mstatus_d_wpri4__57_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__56_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__56_ <= mstatus_d_wpri4__56_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__55_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__55_ <= mstatus_d_wpri4__55_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__54_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__54_ <= mstatus_d_wpri4__54_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__53_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__53_ <= mstatus_d_wpri4__53_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__52_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__52_ <= mstatus_d_wpri4__52_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__51_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__51_ <= mstatus_d_wpri4__51_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__50_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__50_ <= mstatus_d_wpri4__50_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__49_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__49_ <= mstatus_d_wpri4__49_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__48_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__48_ <= mstatus_d_wpri4__48_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__47_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__47_ <= mstatus_d_wpri4__47_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__46_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__46_ <= mstatus_d_wpri4__46_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__45_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__45_ <= mstatus_d_wpri4__45_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__44_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__44_ <= mstatus_d_wpri4__44_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__43_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__43_ <= mstatus_d_wpri4__43_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__42_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__42_ <= mstatus_d_wpri4__42_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__41_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__41_ <= mstatus_d_wpri4__41_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__40_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__40_ <= mstatus_d_wpri4__40_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__39_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__39_ <= mstatus_d_wpri4__39_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__38_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__38_ <= mstatus_d_wpri4__38_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__37_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__37_ <= mstatus_d_wpri4__37_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri4__36_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri4__36_ <= mstatus_d_wpri4__36_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_sxl__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_sxl__1_ <= 1'b1;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_sxl__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_sxl__0_ <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_uxl__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_uxl__1_ <= 1'b1;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_uxl__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_uxl__0_ <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__8_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__8_ <= mstatus_d_wpri3__8_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__7_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__7_ <= mstatus_d_wpri3__7_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__6_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__6_ <= mstatus_d_wpri3__6_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__5_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__5_ <= mstatus_d_wpri3__5_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__4_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__4_ <= mstatus_d_wpri3__4_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__3_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__3_ <= mstatus_d_wpri3__3_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__2_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__2_ <= mstatus_d_wpri3__2_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__1_ <= mstatus_d_wpri3__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri3__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri3__0_ <= mstatus_d_wpri3__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      tsr_o <= 1'b0;
    end else if(1'b1) begin
      tsr_o <= mstatus_d_tsr_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      tw_o <= 1'b0;
    end else if(1'b1) begin
      tw_o <= mstatus_d_tw_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      tvm_o <= 1'b0;
    end else if(1'b1) begin
      tvm_o <= mstatus_d_tvm_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mxr_o <= 1'b0;
    end else if(1'b1) begin
      mxr_o <= mstatus_d_mxr_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sum_o <= 1'b0;
    end else if(1'b1) begin
      sum_o <= mstatus_d_sum_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_mprv_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mprv_ <= mstatus_d_mprv_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_xs__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_xs__1_ <= mstatus_d_xs__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_xs__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_xs__0_ <= mstatus_d_xs__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fs_o[1] <= 1'b0;
    end else if(1'b1) begin
      fs_o[1] <= mstatus_d_fs__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      fs_o[0] <= 1'b0;
    end else if(1'b1) begin
      fs_o[0] <= mstatus_d_fs__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_mpp__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mpp__1_ <= mstatus_d_mpp__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_mpp__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mpp__0_ <= mstatus_d_mpp__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri2__1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri2__1_ <= mstatus_d_wpri2__1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri2__0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri2__0_ <= mstatus_d_wpri2__0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_spp_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_spp_ <= mstatus_d_spp_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_mpie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mpie_ <= mstatus_d_mpie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri1_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri1_ <= mstatus_d_wpri1_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_spie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_spie_ <= mstatus_d_spie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_upie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_upie_ <= mstatus_d_upie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_mie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mie_ <= mstatus_d_mie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_wpri0_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_wpri0_ <= mstatus_d_wpri0_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_sie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_sie_ <= mstatus_d_sie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mstatus_q_uie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_uie_ <= mstatus_d_uie_;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_rst_load_q <= 1'b1;
    end else if(1'b1) begin
      mtvec_rst_load_q <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[63] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[63] <= mtvec_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[62] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[62] <= mtvec_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[61] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[61] <= mtvec_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[60] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[60] <= mtvec_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[59] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[59] <= mtvec_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[58] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[58] <= mtvec_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[57] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[57] <= mtvec_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[56] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[56] <= mtvec_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[55] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[55] <= mtvec_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[54] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[54] <= mtvec_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[53] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[53] <= mtvec_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[52] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[52] <= mtvec_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[51] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[51] <= mtvec_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[50] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[50] <= mtvec_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[49] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[49] <= mtvec_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[48] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[48] <= mtvec_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[47] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[47] <= mtvec_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[46] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[46] <= mtvec_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[45] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[45] <= mtvec_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[44] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[44] <= mtvec_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[43] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[43] <= mtvec_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[42] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[42] <= mtvec_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[41] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[41] <= mtvec_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[40] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[40] <= mtvec_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[39] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[39] <= mtvec_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[38] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[38] <= mtvec_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[37] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[37] <= mtvec_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[36] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[36] <= mtvec_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[35] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[35] <= mtvec_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[34] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[34] <= mtvec_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[33] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[33] <= mtvec_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[32] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[32] <= mtvec_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[31] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[31] <= mtvec_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[30] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[30] <= mtvec_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[29] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[29] <= mtvec_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[28] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[28] <= mtvec_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[27] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[27] <= mtvec_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[26] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[26] <= mtvec_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[25] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[25] <= mtvec_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[24] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[24] <= mtvec_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[23] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[23] <= mtvec_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[22] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[22] <= mtvec_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[21] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[21] <= mtvec_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[20] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[20] <= mtvec_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[19] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[19] <= mtvec_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[18] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[18] <= mtvec_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[17] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[17] <= mtvec_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[16] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[16] <= mtvec_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[15] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[15] <= mtvec_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[14] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[14] <= mtvec_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[13] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[13] <= mtvec_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[12] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[12] <= mtvec_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[11] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[11] <= mtvec_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[10] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[10] <= mtvec_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[9] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[9] <= mtvec_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[8] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[8] <= mtvec_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[7] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[7] <= mtvec_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[6] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[6] <= mtvec_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[5] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[5] <= mtvec_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[4] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[4] <= mtvec_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[3] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[3] <= mtvec_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[2] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[2] <= mtvec_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[1] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[1] <= mtvec_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtvec_q[0] <= 1'b0;
    end else if(1'b1) begin
      mtvec_q[0] <= mtvec_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[63] <= 1'b0;
    end else begin
      medeleg_d[63] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[62] <= 1'b0;
    end else begin
      medeleg_d[62] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[61] <= 1'b0;
    end else begin
      medeleg_d[61] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[60] <= 1'b0;
    end else begin
      medeleg_d[60] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[59] <= 1'b0;
    end else begin
      medeleg_d[59] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[58] <= 1'b0;
    end else begin
      medeleg_d[58] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[57] <= 1'b0;
    end else begin
      medeleg_d[57] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[56] <= 1'b0;
    end else begin
      medeleg_d[56] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[55] <= 1'b0;
    end else begin
      medeleg_d[55] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[54] <= 1'b0;
    end else begin
      medeleg_d[54] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[53] <= 1'b0;
    end else begin
      medeleg_d[53] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[52] <= 1'b0;
    end else begin
      medeleg_d[52] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[51] <= 1'b0;
    end else begin
      medeleg_d[51] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[50] <= 1'b0;
    end else begin
      medeleg_d[50] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[49] <= 1'b0;
    end else begin
      medeleg_d[49] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[48] <= 1'b0;
    end else begin
      medeleg_d[48] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[47] <= 1'b0;
    end else begin
      medeleg_d[47] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[46] <= 1'b0;
    end else begin
      medeleg_d[46] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[45] <= 1'b0;
    end else begin
      medeleg_d[45] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[44] <= 1'b0;
    end else begin
      medeleg_d[44] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[43] <= 1'b0;
    end else begin
      medeleg_d[43] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[42] <= 1'b0;
    end else begin
      medeleg_d[42] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[41] <= 1'b0;
    end else begin
      medeleg_d[41] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[40] <= 1'b0;
    end else begin
      medeleg_d[40] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[39] <= 1'b0;
    end else begin
      medeleg_d[39] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[38] <= 1'b0;
    end else begin
      medeleg_d[38] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[37] <= 1'b0;
    end else begin
      medeleg_d[37] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[36] <= 1'b0;
    end else begin
      medeleg_d[36] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[35] <= 1'b0;
    end else begin
      medeleg_d[35] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[34] <= 1'b0;
    end else begin
      medeleg_d[34] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[33] <= 1'b0;
    end else begin
      medeleg_d[33] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[32] <= 1'b0;
    end else begin
      medeleg_d[32] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[31] <= 1'b0;
    end else begin
      medeleg_d[31] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[30] <= 1'b0;
    end else begin
      medeleg_d[30] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[29] <= 1'b0;
    end else begin
      medeleg_d[29] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[28] <= 1'b0;
    end else begin
      medeleg_d[28] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[27] <= 1'b0;
    end else begin
      medeleg_d[27] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[26] <= 1'b0;
    end else begin
      medeleg_d[26] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[25] <= 1'b0;
    end else begin
      medeleg_d[25] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[24] <= 1'b0;
    end else begin
      medeleg_d[24] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[23] <= 1'b0;
    end else begin
      medeleg_d[23] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[22] <= 1'b0;
    end else begin
      medeleg_d[22] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[21] <= 1'b0;
    end else begin
      medeleg_d[21] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[20] <= 1'b0;
    end else begin
      medeleg_d[20] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[19] <= 1'b0;
    end else begin
      medeleg_d[19] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[18] <= 1'b0;
    end else begin
      medeleg_d[18] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[17] <= 1'b0;
    end else begin
      medeleg_d[17] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[16] <= 1'b0;
    end else begin
      medeleg_d[16] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q_15 <= 1'b0;
    end else if(1'b1) begin
      medeleg_q_15 <= medeleg_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[14] <= 1'b0;
    end else begin
      medeleg_d[14] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q[13] <= 1'b0;
    end else if(1'b1) begin
      medeleg_q[13] <= medeleg_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q[12] <= 1'b0;
    end else if(1'b1) begin
      medeleg_q[12] <= medeleg_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[11] <= 1'b0;
    end else begin
      medeleg_d[11] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[10] <= 1'b0;
    end else begin
      medeleg_d[10] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[9] <= 1'b0;
    end else begin
      medeleg_d[9] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q_8 <= 1'b0;
    end else if(1'b1) begin
      medeleg_q_8 <= medeleg_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[7] <= 1'b0;
    end else begin
      medeleg_d[7] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[6] <= 1'b0;
    end else begin
      medeleg_d[6] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[5] <= 1'b0;
    end else begin
      medeleg_d[5] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[4] <= 1'b0;
    end else begin
      medeleg_d[4] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q_3 <= 1'b0;
    end else if(1'b1) begin
      medeleg_q_3 <= medeleg_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[2] <= 1'b0;
    end else begin
      medeleg_d[2] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_d[1] <= 1'b0;
    end else begin
      medeleg_d[1] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      medeleg_q_0 <= 1'b0;
    end else if(1'b1) begin
      medeleg_q_0 <= medeleg_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[63] <= 1'b0;
    end else begin
      mideleg_d[63] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[62] <= 1'b0;
    end else begin
      mideleg_d[62] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[61] <= 1'b0;
    end else begin
      mideleg_d[61] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[60] <= 1'b0;
    end else begin
      mideleg_d[60] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[59] <= 1'b0;
    end else begin
      mideleg_d[59] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[58] <= 1'b0;
    end else begin
      mideleg_d[58] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[57] <= 1'b0;
    end else begin
      mideleg_d[57] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[56] <= 1'b0;
    end else begin
      mideleg_d[56] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[55] <= 1'b0;
    end else begin
      mideleg_d[55] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[54] <= 1'b0;
    end else begin
      mideleg_d[54] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[53] <= 1'b0;
    end else begin
      mideleg_d[53] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[52] <= 1'b0;
    end else begin
      mideleg_d[52] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[51] <= 1'b0;
    end else begin
      mideleg_d[51] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[50] <= 1'b0;
    end else begin
      mideleg_d[50] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[49] <= 1'b0;
    end else begin
      mideleg_d[49] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[48] <= 1'b0;
    end else begin
      mideleg_d[48] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[47] <= 1'b0;
    end else begin
      mideleg_d[47] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[46] <= 1'b0;
    end else begin
      mideleg_d[46] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[45] <= 1'b0;
    end else begin
      mideleg_d[45] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[44] <= 1'b0;
    end else begin
      mideleg_d[44] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[43] <= 1'b0;
    end else begin
      mideleg_d[43] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[42] <= 1'b0;
    end else begin
      mideleg_d[42] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[41] <= 1'b0;
    end else begin
      mideleg_d[41] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[40] <= 1'b0;
    end else begin
      mideleg_d[40] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[39] <= 1'b0;
    end else begin
      mideleg_d[39] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[38] <= 1'b0;
    end else begin
      mideleg_d[38] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[37] <= 1'b0;
    end else begin
      mideleg_d[37] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[36] <= 1'b0;
    end else begin
      mideleg_d[36] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[35] <= 1'b0;
    end else begin
      mideleg_d[35] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[34] <= 1'b0;
    end else begin
      mideleg_d[34] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[33] <= 1'b0;
    end else begin
      mideleg_d[33] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[32] <= 1'b0;
    end else begin
      mideleg_d[32] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[31] <= 1'b0;
    end else begin
      mideleg_d[31] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[30] <= 1'b0;
    end else begin
      mideleg_d[30] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[29] <= 1'b0;
    end else begin
      mideleg_d[29] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[28] <= 1'b0;
    end else begin
      mideleg_d[28] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[27] <= 1'b0;
    end else begin
      mideleg_d[27] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[26] <= 1'b0;
    end else begin
      mideleg_d[26] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[25] <= 1'b0;
    end else begin
      mideleg_d[25] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[24] <= 1'b0;
    end else begin
      mideleg_d[24] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[23] <= 1'b0;
    end else begin
      mideleg_d[23] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[22] <= 1'b0;
    end else begin
      mideleg_d[22] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[21] <= 1'b0;
    end else begin
      mideleg_d[21] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[20] <= 1'b0;
    end else begin
      mideleg_d[20] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[19] <= 1'b0;
    end else begin
      mideleg_d[19] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[18] <= 1'b0;
    end else begin
      mideleg_d[18] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[17] <= 1'b0;
    end else begin
      mideleg_d[17] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[16] <= 1'b0;
    end else begin
      mideleg_d[16] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[15] <= 1'b0;
    end else begin
      mideleg_d[15] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[14] <= 1'b0;
    end else begin
      mideleg_d[14] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[13] <= 1'b0;
    end else begin
      mideleg_d[13] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[12] <= 1'b0;
    end else begin
      mideleg_d[12] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[11] <= 1'b0;
    end else begin
      mideleg_d[11] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[10] <= 1'b0;
    end else begin
      mideleg_d[10] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_q[9] <= 1'b0;
    end else if(1'b1) begin
      mideleg_q[9] <= mideleg_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[8] <= 1'b0;
    end else begin
      mideleg_d[8] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[7] <= 1'b0;
    end else begin
      mideleg_d[7] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[6] <= 1'b0;
    end else begin
      mideleg_d[6] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_q_5 <= 1'b0;
    end else if(1'b1) begin
      mideleg_q_5 <= mideleg_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[4] <= 1'b0;
    end else begin
      mideleg_d[4] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[3] <= 1'b0;
    end else begin
      mideleg_d[3] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[2] <= 1'b0;
    end else begin
      mideleg_d[2] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_q_1 <= 1'b0;
    end else if(1'b1) begin
      mideleg_q_1 <= mideleg_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mideleg_d[0] <= 1'b0;
    end else begin
      mideleg_d[0] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[63] <= 1'b0;
    end else begin
      mip_d[63] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[62] <= 1'b0;
    end else begin
      mip_d[62] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[61] <= 1'b0;
    end else begin
      mip_d[61] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[60] <= 1'b0;
    end else begin
      mip_d[60] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[59] <= 1'b0;
    end else begin
      mip_d[59] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[58] <= 1'b0;
    end else begin
      mip_d[58] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[57] <= 1'b0;
    end else begin
      mip_d[57] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[56] <= 1'b0;
    end else begin
      mip_d[56] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[55] <= 1'b0;
    end else begin
      mip_d[55] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[54] <= 1'b0;
    end else begin
      mip_d[54] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[53] <= 1'b0;
    end else begin
      mip_d[53] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[52] <= 1'b0;
    end else begin
      mip_d[52] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[51] <= 1'b0;
    end else begin
      mip_d[51] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[50] <= 1'b0;
    end else begin
      mip_d[50] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[49] <= 1'b0;
    end else begin
      mip_d[49] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[48] <= 1'b0;
    end else begin
      mip_d[48] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[47] <= 1'b0;
    end else begin
      mip_d[47] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[46] <= 1'b0;
    end else begin
      mip_d[46] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[45] <= 1'b0;
    end else begin
      mip_d[45] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[44] <= 1'b0;
    end else begin
      mip_d[44] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[43] <= 1'b0;
    end else begin
      mip_d[43] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[42] <= 1'b0;
    end else begin
      mip_d[42] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[41] <= 1'b0;
    end else begin
      mip_d[41] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[40] <= 1'b0;
    end else begin
      mip_d[40] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[39] <= 1'b0;
    end else begin
      mip_d[39] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[38] <= 1'b0;
    end else begin
      mip_d[38] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[37] <= 1'b0;
    end else begin
      mip_d[37] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[36] <= 1'b0;
    end else begin
      mip_d[36] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[35] <= 1'b0;
    end else begin
      mip_d[35] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[34] <= 1'b0;
    end else begin
      mip_d[34] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[33] <= 1'b0;
    end else begin
      mip_d[33] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[32] <= 1'b0;
    end else begin
      mip_d[32] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[31] <= 1'b0;
    end else begin
      mip_d[31] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[30] <= 1'b0;
    end else begin
      mip_d[30] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[29] <= 1'b0;
    end else begin
      mip_d[29] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[28] <= 1'b0;
    end else begin
      mip_d[28] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[27] <= 1'b0;
    end else begin
      mip_d[27] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[26] <= 1'b0;
    end else begin
      mip_d[26] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[25] <= 1'b0;
    end else begin
      mip_d[25] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[24] <= 1'b0;
    end else begin
      mip_d[24] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[23] <= 1'b0;
    end else begin
      mip_d[23] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[22] <= 1'b0;
    end else begin
      mip_d[22] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[21] <= 1'b0;
    end else begin
      mip_d[21] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[20] <= 1'b0;
    end else begin
      mip_d[20] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[19] <= 1'b0;
    end else begin
      mip_d[19] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[18] <= 1'b0;
    end else begin
      mip_d[18] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[17] <= 1'b0;
    end else begin
      mip_d[17] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[16] <= 1'b0;
    end else begin
      mip_d[16] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[15] <= 1'b0;
    end else begin
      mip_d[15] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[14] <= 1'b0;
    end else begin
      mip_d[14] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[13] <= 1'b0;
    end else begin
      mip_d[13] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d[12] <= 1'b0;
    end else begin
      mip_d[12] <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q[11] <= 1'b0;
    end else if(1'b1) begin
      mip_q[11] <= irq_i[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_10 <= 1'b0;
    end else begin
      mip_d_10 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q_9 <= 1'b0;
    end else if(1'b1) begin
      mip_q_9 <= mip_d_9;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_8 <= 1'b0;
    end else begin
      mip_d_8 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q_7 <= 1'b0;
    end else if(1'b1) begin
      mip_q_7 <= time_irq_i;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_6 <= 1'b0;
    end else begin
      mip_d_6 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q_5 <= 1'b0;
    end else if(1'b1) begin
      mip_q_5 <= mip_d_5;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_4 <= 1'b0;
    end else begin
      mip_d_4 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q_3 <= 1'b0;
    end else if(1'b1) begin
      mip_q_3 <= ipi_i;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_2 <= 1'b0;
    end else begin
      mip_d_2 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_q_1 <= 1'b0;
    end else if(1'b1) begin
      mip_q_1 <= mip_d_1;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mip_d_0 <= 1'b0;
    end else begin
      mip_d_0 <= N168;
    end
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[63] <= 1'b0;
    end else if(1'b1) begin
      mie_q[63] <= mie_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[62] <= 1'b0;
    end else if(1'b1) begin
      mie_q[62] <= mie_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[61] <= 1'b0;
    end else if(1'b1) begin
      mie_q[61] <= mie_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[60] <= 1'b0;
    end else if(1'b1) begin
      mie_q[60] <= mie_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[59] <= 1'b0;
    end else if(1'b1) begin
      mie_q[59] <= mie_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[58] <= 1'b0;
    end else if(1'b1) begin
      mie_q[58] <= mie_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[57] <= 1'b0;
    end else if(1'b1) begin
      mie_q[57] <= mie_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[56] <= 1'b0;
    end else if(1'b1) begin
      mie_q[56] <= mie_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[55] <= 1'b0;
    end else if(1'b1) begin
      mie_q[55] <= mie_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[54] <= 1'b0;
    end else if(1'b1) begin
      mie_q[54] <= mie_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[53] <= 1'b0;
    end else if(1'b1) begin
      mie_q[53] <= mie_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[52] <= 1'b0;
    end else if(1'b1) begin
      mie_q[52] <= mie_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[51] <= 1'b0;
    end else if(1'b1) begin
      mie_q[51] <= mie_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[50] <= 1'b0;
    end else if(1'b1) begin
      mie_q[50] <= mie_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[49] <= 1'b0;
    end else if(1'b1) begin
      mie_q[49] <= mie_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[48] <= 1'b0;
    end else if(1'b1) begin
      mie_q[48] <= mie_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[47] <= 1'b0;
    end else if(1'b1) begin
      mie_q[47] <= mie_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[46] <= 1'b0;
    end else if(1'b1) begin
      mie_q[46] <= mie_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[45] <= 1'b0;
    end else if(1'b1) begin
      mie_q[45] <= mie_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[44] <= 1'b0;
    end else if(1'b1) begin
      mie_q[44] <= mie_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[43] <= 1'b0;
    end else if(1'b1) begin
      mie_q[43] <= mie_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[42] <= 1'b0;
    end else if(1'b1) begin
      mie_q[42] <= mie_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[41] <= 1'b0;
    end else if(1'b1) begin
      mie_q[41] <= mie_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[40] <= 1'b0;
    end else if(1'b1) begin
      mie_q[40] <= mie_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[39] <= 1'b0;
    end else if(1'b1) begin
      mie_q[39] <= mie_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[38] <= 1'b0;
    end else if(1'b1) begin
      mie_q[38] <= mie_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[37] <= 1'b0;
    end else if(1'b1) begin
      mie_q[37] <= mie_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[36] <= 1'b0;
    end else if(1'b1) begin
      mie_q[36] <= mie_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[35] <= 1'b0;
    end else if(1'b1) begin
      mie_q[35] <= mie_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[34] <= 1'b0;
    end else if(1'b1) begin
      mie_q[34] <= mie_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[33] <= 1'b0;
    end else if(1'b1) begin
      mie_q[33] <= mie_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[32] <= 1'b0;
    end else if(1'b1) begin
      mie_q[32] <= mie_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[31] <= 1'b0;
    end else if(1'b1) begin
      mie_q[31] <= mie_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[30] <= 1'b0;
    end else if(1'b1) begin
      mie_q[30] <= mie_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[29] <= 1'b0;
    end else if(1'b1) begin
      mie_q[29] <= mie_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[28] <= 1'b0;
    end else if(1'b1) begin
      mie_q[28] <= mie_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[27] <= 1'b0;
    end else if(1'b1) begin
      mie_q[27] <= mie_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[26] <= 1'b0;
    end else if(1'b1) begin
      mie_q[26] <= mie_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[25] <= 1'b0;
    end else if(1'b1) begin
      mie_q[25] <= mie_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[24] <= 1'b0;
    end else if(1'b1) begin
      mie_q[24] <= mie_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[23] <= 1'b0;
    end else if(1'b1) begin
      mie_q[23] <= mie_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[22] <= 1'b0;
    end else if(1'b1) begin
      mie_q[22] <= mie_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[21] <= 1'b0;
    end else if(1'b1) begin
      mie_q[21] <= mie_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[20] <= 1'b0;
    end else if(1'b1) begin
      mie_q[20] <= mie_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[19] <= 1'b0;
    end else if(1'b1) begin
      mie_q[19] <= mie_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[18] <= 1'b0;
    end else if(1'b1) begin
      mie_q[18] <= mie_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[17] <= 1'b0;
    end else if(1'b1) begin
      mie_q[17] <= mie_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[16] <= 1'b0;
    end else if(1'b1) begin
      mie_q[16] <= mie_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[15] <= 1'b0;
    end else if(1'b1) begin
      mie_q[15] <= mie_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[14] <= 1'b0;
    end else if(1'b1) begin
      mie_q[14] <= mie_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[13] <= 1'b0;
    end else if(1'b1) begin
      mie_q[13] <= mie_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[12] <= 1'b0;
    end else if(1'b1) begin
      mie_q[12] <= mie_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[11] <= 1'b0;
    end else if(1'b1) begin
      mie_q[11] <= mie_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[10] <= 1'b0;
    end else if(1'b1) begin
      mie_q[10] <= mie_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[9] <= 1'b0;
    end else if(1'b1) begin
      mie_q[9] <= mie_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[8] <= 1'b0;
    end else if(1'b1) begin
      mie_q[8] <= mie_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[7] <= 1'b0;
    end else if(1'b1) begin
      mie_q[7] <= mie_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[6] <= 1'b0;
    end else if(1'b1) begin
      mie_q[6] <= mie_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[5] <= 1'b0;
    end else if(1'b1) begin
      mie_q[5] <= mie_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[4] <= 1'b0;
    end else if(1'b1) begin
      mie_q[4] <= mie_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[3] <= 1'b0;
    end else if(1'b1) begin
      mie_q[3] <= mie_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[2] <= 1'b0;
    end else if(1'b1) begin
      mie_q[2] <= mie_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[1] <= 1'b0;
    end else if(1'b1) begin
      mie_q[1] <= mie_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mie_q[0] <= 1'b0;
    end else if(1'b1) begin
      mie_q[0] <= mie_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[63] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[63] <= mepc_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[62] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[62] <= mepc_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[61] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[61] <= mepc_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[60] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[60] <= mepc_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[59] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[59] <= mepc_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[58] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[58] <= mepc_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[57] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[57] <= mepc_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[56] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[56] <= mepc_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[55] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[55] <= mepc_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[54] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[54] <= mepc_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[53] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[53] <= mepc_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[52] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[52] <= mepc_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[51] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[51] <= mepc_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[50] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[50] <= mepc_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[49] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[49] <= mepc_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[48] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[48] <= mepc_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[47] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[47] <= mepc_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[46] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[46] <= mepc_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[45] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[45] <= mepc_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[44] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[44] <= mepc_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[43] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[43] <= mepc_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[42] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[42] <= mepc_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[41] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[41] <= mepc_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[40] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[40] <= mepc_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[39] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[39] <= mepc_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[38] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[38] <= mepc_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[37] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[37] <= mepc_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[36] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[36] <= mepc_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[35] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[35] <= mepc_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[34] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[34] <= mepc_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[33] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[33] <= mepc_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[32] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[32] <= mepc_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[31] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[31] <= mepc_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[30] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[30] <= mepc_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[29] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[29] <= mepc_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[28] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[28] <= mepc_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[27] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[27] <= mepc_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[26] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[26] <= mepc_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[25] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[25] <= mepc_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[24] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[24] <= mepc_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[23] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[23] <= mepc_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[22] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[22] <= mepc_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[21] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[21] <= mepc_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[20] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[20] <= mepc_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[19] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[19] <= mepc_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[18] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[18] <= mepc_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[17] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[17] <= mepc_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[16] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[16] <= mepc_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[15] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[15] <= mepc_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[14] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[14] <= mepc_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[13] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[13] <= mepc_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[12] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[12] <= mepc_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[11] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[11] <= mepc_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[10] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[10] <= mepc_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[9] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[9] <= mepc_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[8] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[8] <= mepc_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[7] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[7] <= mepc_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[6] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[6] <= mepc_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[5] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[5] <= mepc_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[4] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[4] <= mepc_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[3] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[3] <= mepc_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[2] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[2] <= mepc_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[1] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[1] <= mepc_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mepc_q[0] <= 1'b0;
    end else if(1'b1) begin
      mepc_q[0] <= mepc_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[63] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[63] <= mcause_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[62] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[62] <= mcause_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[61] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[61] <= mcause_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[60] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[60] <= mcause_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[59] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[59] <= mcause_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[58] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[58] <= mcause_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[57] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[57] <= mcause_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[56] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[56] <= mcause_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[55] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[55] <= mcause_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[54] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[54] <= mcause_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[53] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[53] <= mcause_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[52] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[52] <= mcause_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[51] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[51] <= mcause_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[50] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[50] <= mcause_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[49] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[49] <= mcause_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[48] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[48] <= mcause_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[47] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[47] <= mcause_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[46] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[46] <= mcause_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[45] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[45] <= mcause_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[44] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[44] <= mcause_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[43] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[43] <= mcause_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[42] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[42] <= mcause_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[41] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[41] <= mcause_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[40] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[40] <= mcause_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[39] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[39] <= mcause_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[38] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[38] <= mcause_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[37] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[37] <= mcause_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[36] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[36] <= mcause_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[35] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[35] <= mcause_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[34] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[34] <= mcause_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[33] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[33] <= mcause_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[32] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[32] <= mcause_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[31] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[31] <= mcause_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[30] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[30] <= mcause_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[29] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[29] <= mcause_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[28] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[28] <= mcause_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[27] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[27] <= mcause_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[26] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[26] <= mcause_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[25] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[25] <= mcause_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[24] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[24] <= mcause_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[23] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[23] <= mcause_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[22] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[22] <= mcause_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[21] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[21] <= mcause_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[20] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[20] <= mcause_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[19] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[19] <= mcause_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[18] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[18] <= mcause_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[17] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[17] <= mcause_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[16] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[16] <= mcause_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[15] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[15] <= mcause_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[14] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[14] <= mcause_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[13] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[13] <= mcause_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[12] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[12] <= mcause_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[11] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[11] <= mcause_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[10] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[10] <= mcause_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[9] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[9] <= mcause_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[8] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[8] <= mcause_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[7] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[7] <= mcause_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[6] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[6] <= mcause_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[5] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[5] <= mcause_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[4] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[4] <= mcause_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[3] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[3] <= mcause_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[2] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[2] <= mcause_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[1] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[1] <= mcause_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mcause_q[0] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[0] <= mcause_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[63] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[63] <= mscratch_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[62] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[62] <= mscratch_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[61] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[61] <= mscratch_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[60] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[60] <= mscratch_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[59] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[59] <= mscratch_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[58] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[58] <= mscratch_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[57] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[57] <= mscratch_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[56] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[56] <= mscratch_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[55] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[55] <= mscratch_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[54] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[54] <= mscratch_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[53] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[53] <= mscratch_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[52] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[52] <= mscratch_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[51] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[51] <= mscratch_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[50] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[50] <= mscratch_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[49] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[49] <= mscratch_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[48] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[48] <= mscratch_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[47] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[47] <= mscratch_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[46] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[46] <= mscratch_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[45] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[45] <= mscratch_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[44] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[44] <= mscratch_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[43] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[43] <= mscratch_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[42] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[42] <= mscratch_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[41] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[41] <= mscratch_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[40] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[40] <= mscratch_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[39] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[39] <= mscratch_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[38] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[38] <= mscratch_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[37] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[37] <= mscratch_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[36] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[36] <= mscratch_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[35] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[35] <= mscratch_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[34] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[34] <= mscratch_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[33] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[33] <= mscratch_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[32] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[32] <= mscratch_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[31] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[31] <= mscratch_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[30] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[30] <= mscratch_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[29] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[29] <= mscratch_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[28] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[28] <= mscratch_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[27] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[27] <= mscratch_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[26] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[26] <= mscratch_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[25] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[25] <= mscratch_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[24] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[24] <= mscratch_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[23] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[23] <= mscratch_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[22] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[22] <= mscratch_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[21] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[21] <= mscratch_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[20] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[20] <= mscratch_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[19] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[19] <= mscratch_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[18] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[18] <= mscratch_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[17] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[17] <= mscratch_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[16] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[16] <= mscratch_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[15] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[15] <= mscratch_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[14] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[14] <= mscratch_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[13] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[13] <= mscratch_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[12] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[12] <= mscratch_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[11] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[11] <= mscratch_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[10] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[10] <= mscratch_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[9] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[9] <= mscratch_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[8] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[8] <= mscratch_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[7] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[7] <= mscratch_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[6] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[6] <= mscratch_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[5] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[5] <= mscratch_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[4] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[4] <= mscratch_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[3] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[3] <= mscratch_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[2] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[2] <= mscratch_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[1] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[1] <= mscratch_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mscratch_q[0] <= 1'b0;
    end else if(1'b1) begin
      mscratch_q[0] <= mscratch_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[63] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[63] <= mtval_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[62] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[62] <= mtval_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[61] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[61] <= mtval_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[60] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[60] <= mtval_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[59] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[59] <= mtval_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[58] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[58] <= mtval_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[57] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[57] <= mtval_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[56] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[56] <= mtval_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[55] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[55] <= mtval_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[54] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[54] <= mtval_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[53] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[53] <= mtval_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[52] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[52] <= mtval_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[51] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[51] <= mtval_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[50] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[50] <= mtval_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[49] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[49] <= mtval_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[48] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[48] <= mtval_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[47] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[47] <= mtval_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[46] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[46] <= mtval_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[45] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[45] <= mtval_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[44] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[44] <= mtval_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[43] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[43] <= mtval_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[42] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[42] <= mtval_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[41] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[41] <= mtval_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[40] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[40] <= mtval_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[39] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[39] <= mtval_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[38] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[38] <= mtval_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[37] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[37] <= mtval_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[36] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[36] <= mtval_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[35] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[35] <= mtval_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[34] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[34] <= mtval_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[33] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[33] <= mtval_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[32] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[32] <= mtval_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[31] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[31] <= mtval_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[30] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[30] <= mtval_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[29] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[29] <= mtval_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[28] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[28] <= mtval_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[27] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[27] <= mtval_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[26] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[26] <= mtval_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[25] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[25] <= mtval_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[24] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[24] <= mtval_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[23] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[23] <= mtval_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[22] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[22] <= mtval_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[21] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[21] <= mtval_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[20] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[20] <= mtval_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[19] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[19] <= mtval_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[18] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[18] <= mtval_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[17] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[17] <= mtval_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[16] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[16] <= mtval_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[15] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[15] <= mtval_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[14] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[14] <= mtval_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[13] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[13] <= mtval_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[12] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[12] <= mtval_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[11] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[11] <= mtval_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[10] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[10] <= mtval_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[9] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[9] <= mtval_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[8] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[8] <= mtval_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[7] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[7] <= mtval_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[6] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[6] <= mtval_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[5] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[5] <= mtval_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[4] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[4] <= mtval_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[3] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[3] <= mtval_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[2] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[2] <= mtval_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[1] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[1] <= mtval_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      mtval_q[0] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[0] <= mtval_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[63] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[63] <= dcache_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[62] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[62] <= dcache_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[61] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[61] <= dcache_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[60] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[60] <= dcache_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[59] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[59] <= dcache_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[58] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[58] <= dcache_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[57] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[57] <= dcache_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[56] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[56] <= dcache_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[55] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[55] <= dcache_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[54] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[54] <= dcache_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[53] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[53] <= dcache_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[52] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[52] <= dcache_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[51] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[51] <= dcache_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[50] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[50] <= dcache_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[49] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[49] <= dcache_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[48] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[48] <= dcache_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[47] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[47] <= dcache_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[46] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[46] <= dcache_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[45] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[45] <= dcache_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[44] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[44] <= dcache_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[43] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[43] <= dcache_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[42] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[42] <= dcache_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[41] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[41] <= dcache_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[40] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[40] <= dcache_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[39] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[39] <= dcache_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[38] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[38] <= dcache_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[37] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[37] <= dcache_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[36] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[36] <= dcache_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[35] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[35] <= dcache_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[34] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[34] <= dcache_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[33] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[33] <= dcache_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[32] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[32] <= dcache_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[31] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[31] <= dcache_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[30] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[30] <= dcache_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[29] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[29] <= dcache_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[28] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[28] <= dcache_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[27] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[27] <= dcache_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[26] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[26] <= dcache_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[25] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[25] <= dcache_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[24] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[24] <= dcache_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[23] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[23] <= dcache_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[22] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[22] <= dcache_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[21] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[21] <= dcache_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[20] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[20] <= dcache_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[19] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[19] <= dcache_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[18] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[18] <= dcache_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[17] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[17] <= dcache_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[16] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[16] <= dcache_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[15] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[15] <= dcache_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[14] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[14] <= dcache_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[13] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[13] <= dcache_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[12] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[12] <= dcache_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[11] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[11] <= dcache_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[10] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[10] <= dcache_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[9] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[9] <= dcache_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[8] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[8] <= dcache_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[7] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[7] <= dcache_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[6] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[6] <= dcache_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[5] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[5] <= dcache_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[4] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[4] <= dcache_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[3] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[3] <= dcache_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[2] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[2] <= dcache_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_q[1] <= 1'b0;
    end else if(1'b1) begin
      dcache_q[1] <= dcache_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      dcache_en_o <= 1'b1;
    end else if(1'b1) begin
      dcache_en_o <= dcache_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[63] <= 1'b0;
    end else if(1'b1) begin
      icache_q[63] <= icache_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[62] <= 1'b0;
    end else if(1'b1) begin
      icache_q[62] <= icache_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[61] <= 1'b0;
    end else if(1'b1) begin
      icache_q[61] <= icache_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[60] <= 1'b0;
    end else if(1'b1) begin
      icache_q[60] <= icache_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[59] <= 1'b0;
    end else if(1'b1) begin
      icache_q[59] <= icache_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[58] <= 1'b0;
    end else if(1'b1) begin
      icache_q[58] <= icache_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[57] <= 1'b0;
    end else if(1'b1) begin
      icache_q[57] <= icache_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[56] <= 1'b0;
    end else if(1'b1) begin
      icache_q[56] <= icache_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[55] <= 1'b0;
    end else if(1'b1) begin
      icache_q[55] <= icache_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[54] <= 1'b0;
    end else if(1'b1) begin
      icache_q[54] <= icache_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[53] <= 1'b0;
    end else if(1'b1) begin
      icache_q[53] <= icache_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[52] <= 1'b0;
    end else if(1'b1) begin
      icache_q[52] <= icache_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[51] <= 1'b0;
    end else if(1'b1) begin
      icache_q[51] <= icache_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[50] <= 1'b0;
    end else if(1'b1) begin
      icache_q[50] <= icache_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[49] <= 1'b0;
    end else if(1'b1) begin
      icache_q[49] <= icache_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[48] <= 1'b0;
    end else if(1'b1) begin
      icache_q[48] <= icache_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[47] <= 1'b0;
    end else if(1'b1) begin
      icache_q[47] <= icache_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[46] <= 1'b0;
    end else if(1'b1) begin
      icache_q[46] <= icache_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[45] <= 1'b0;
    end else if(1'b1) begin
      icache_q[45] <= icache_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[44] <= 1'b0;
    end else if(1'b1) begin
      icache_q[44] <= icache_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[43] <= 1'b0;
    end else if(1'b1) begin
      icache_q[43] <= icache_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[42] <= 1'b0;
    end else if(1'b1) begin
      icache_q[42] <= icache_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[41] <= 1'b0;
    end else if(1'b1) begin
      icache_q[41] <= icache_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[40] <= 1'b0;
    end else if(1'b1) begin
      icache_q[40] <= icache_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[39] <= 1'b0;
    end else if(1'b1) begin
      icache_q[39] <= icache_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[38] <= 1'b0;
    end else if(1'b1) begin
      icache_q[38] <= icache_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[37] <= 1'b0;
    end else if(1'b1) begin
      icache_q[37] <= icache_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[36] <= 1'b0;
    end else if(1'b1) begin
      icache_q[36] <= icache_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[35] <= 1'b0;
    end else if(1'b1) begin
      icache_q[35] <= icache_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[34] <= 1'b0;
    end else if(1'b1) begin
      icache_q[34] <= icache_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[33] <= 1'b0;
    end else if(1'b1) begin
      icache_q[33] <= icache_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[32] <= 1'b0;
    end else if(1'b1) begin
      icache_q[32] <= icache_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[31] <= 1'b0;
    end else if(1'b1) begin
      icache_q[31] <= icache_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[30] <= 1'b0;
    end else if(1'b1) begin
      icache_q[30] <= icache_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[29] <= 1'b0;
    end else if(1'b1) begin
      icache_q[29] <= icache_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[28] <= 1'b0;
    end else if(1'b1) begin
      icache_q[28] <= icache_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[27] <= 1'b0;
    end else if(1'b1) begin
      icache_q[27] <= icache_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[26] <= 1'b0;
    end else if(1'b1) begin
      icache_q[26] <= icache_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[25] <= 1'b0;
    end else if(1'b1) begin
      icache_q[25] <= icache_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[24] <= 1'b0;
    end else if(1'b1) begin
      icache_q[24] <= icache_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[23] <= 1'b0;
    end else if(1'b1) begin
      icache_q[23] <= icache_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[22] <= 1'b0;
    end else if(1'b1) begin
      icache_q[22] <= icache_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[21] <= 1'b0;
    end else if(1'b1) begin
      icache_q[21] <= icache_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[20] <= 1'b0;
    end else if(1'b1) begin
      icache_q[20] <= icache_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[19] <= 1'b0;
    end else if(1'b1) begin
      icache_q[19] <= icache_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[18] <= 1'b0;
    end else if(1'b1) begin
      icache_q[18] <= icache_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[17] <= 1'b0;
    end else if(1'b1) begin
      icache_q[17] <= icache_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[16] <= 1'b0;
    end else if(1'b1) begin
      icache_q[16] <= icache_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[15] <= 1'b0;
    end else if(1'b1) begin
      icache_q[15] <= icache_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[14] <= 1'b0;
    end else if(1'b1) begin
      icache_q[14] <= icache_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[13] <= 1'b0;
    end else if(1'b1) begin
      icache_q[13] <= icache_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[12] <= 1'b0;
    end else if(1'b1) begin
      icache_q[12] <= icache_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[11] <= 1'b0;
    end else if(1'b1) begin
      icache_q[11] <= icache_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[10] <= 1'b0;
    end else if(1'b1) begin
      icache_q[10] <= icache_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[9] <= 1'b0;
    end else if(1'b1) begin
      icache_q[9] <= icache_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[8] <= 1'b0;
    end else if(1'b1) begin
      icache_q[8] <= icache_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[7] <= 1'b0;
    end else if(1'b1) begin
      icache_q[7] <= icache_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[6] <= 1'b0;
    end else if(1'b1) begin
      icache_q[6] <= icache_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[5] <= 1'b0;
    end else if(1'b1) begin
      icache_q[5] <= icache_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[4] <= 1'b0;
    end else if(1'b1) begin
      icache_q[4] <= icache_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[3] <= 1'b0;
    end else if(1'b1) begin
      icache_q[3] <= icache_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[2] <= 1'b0;
    end else if(1'b1) begin
      icache_q[2] <= icache_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[1] <= 1'b0;
    end else if(1'b1) begin
      icache_q[1] <= icache_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      icache_q[0] <= 1'b1;
    end else if(1'b1) begin
      icache_q[0] <= icache_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[63] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[63] <= sepc_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[62] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[62] <= sepc_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[61] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[61] <= sepc_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[60] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[60] <= sepc_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[59] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[59] <= sepc_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[58] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[58] <= sepc_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[57] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[57] <= sepc_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[56] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[56] <= sepc_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[55] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[55] <= sepc_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[54] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[54] <= sepc_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[53] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[53] <= sepc_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[52] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[52] <= sepc_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[51] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[51] <= sepc_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[50] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[50] <= sepc_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[49] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[49] <= sepc_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[48] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[48] <= sepc_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[47] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[47] <= sepc_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[46] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[46] <= sepc_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[45] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[45] <= sepc_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[44] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[44] <= sepc_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[43] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[43] <= sepc_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[42] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[42] <= sepc_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[41] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[41] <= sepc_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[40] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[40] <= sepc_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[39] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[39] <= sepc_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[38] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[38] <= sepc_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[37] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[37] <= sepc_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[36] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[36] <= sepc_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[35] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[35] <= sepc_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[34] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[34] <= sepc_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[33] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[33] <= sepc_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[32] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[32] <= sepc_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[31] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[31] <= sepc_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[30] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[30] <= sepc_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[29] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[29] <= sepc_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[28] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[28] <= sepc_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[27] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[27] <= sepc_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[26] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[26] <= sepc_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[25] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[25] <= sepc_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[24] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[24] <= sepc_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[23] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[23] <= sepc_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[22] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[22] <= sepc_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[21] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[21] <= sepc_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[20] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[20] <= sepc_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[19] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[19] <= sepc_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[18] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[18] <= sepc_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[17] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[17] <= sepc_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[16] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[16] <= sepc_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[15] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[15] <= sepc_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[14] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[14] <= sepc_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[13] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[13] <= sepc_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[12] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[12] <= sepc_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[11] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[11] <= sepc_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[10] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[10] <= sepc_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[9] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[9] <= sepc_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[8] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[8] <= sepc_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[7] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[7] <= sepc_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[6] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[6] <= sepc_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[5] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[5] <= sepc_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[4] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[4] <= sepc_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[3] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[3] <= sepc_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[2] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[2] <= sepc_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[1] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[1] <= sepc_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sepc_q[0] <= 1'b0;
    end else if(1'b1) begin
      sepc_q[0] <= sepc_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[63] <= 1'b0;
    end else if(1'b1) begin
      scause_q[63] <= scause_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[62] <= 1'b0;
    end else if(1'b1) begin
      scause_q[62] <= scause_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[61] <= 1'b0;
    end else if(1'b1) begin
      scause_q[61] <= scause_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[60] <= 1'b0;
    end else if(1'b1) begin
      scause_q[60] <= scause_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[59] <= 1'b0;
    end else if(1'b1) begin
      scause_q[59] <= scause_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[58] <= 1'b0;
    end else if(1'b1) begin
      scause_q[58] <= scause_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[57] <= 1'b0;
    end else if(1'b1) begin
      scause_q[57] <= scause_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[56] <= 1'b0;
    end else if(1'b1) begin
      scause_q[56] <= scause_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[55] <= 1'b0;
    end else if(1'b1) begin
      scause_q[55] <= scause_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[54] <= 1'b0;
    end else if(1'b1) begin
      scause_q[54] <= scause_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[53] <= 1'b0;
    end else if(1'b1) begin
      scause_q[53] <= scause_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[52] <= 1'b0;
    end else if(1'b1) begin
      scause_q[52] <= scause_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[51] <= 1'b0;
    end else if(1'b1) begin
      scause_q[51] <= scause_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[50] <= 1'b0;
    end else if(1'b1) begin
      scause_q[50] <= scause_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[49] <= 1'b0;
    end else if(1'b1) begin
      scause_q[49] <= scause_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[48] <= 1'b0;
    end else if(1'b1) begin
      scause_q[48] <= scause_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[47] <= 1'b0;
    end else if(1'b1) begin
      scause_q[47] <= scause_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[46] <= 1'b0;
    end else if(1'b1) begin
      scause_q[46] <= scause_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[45] <= 1'b0;
    end else if(1'b1) begin
      scause_q[45] <= scause_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[44] <= 1'b0;
    end else if(1'b1) begin
      scause_q[44] <= scause_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[43] <= 1'b0;
    end else if(1'b1) begin
      scause_q[43] <= scause_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[42] <= 1'b0;
    end else if(1'b1) begin
      scause_q[42] <= scause_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[41] <= 1'b0;
    end else if(1'b1) begin
      scause_q[41] <= scause_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[40] <= 1'b0;
    end else if(1'b1) begin
      scause_q[40] <= scause_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[39] <= 1'b0;
    end else if(1'b1) begin
      scause_q[39] <= scause_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[38] <= 1'b0;
    end else if(1'b1) begin
      scause_q[38] <= scause_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[37] <= 1'b0;
    end else if(1'b1) begin
      scause_q[37] <= scause_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[36] <= 1'b0;
    end else if(1'b1) begin
      scause_q[36] <= scause_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[35] <= 1'b0;
    end else if(1'b1) begin
      scause_q[35] <= scause_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[34] <= 1'b0;
    end else if(1'b1) begin
      scause_q[34] <= scause_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[33] <= 1'b0;
    end else if(1'b1) begin
      scause_q[33] <= scause_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[32] <= 1'b0;
    end else if(1'b1) begin
      scause_q[32] <= scause_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[31] <= 1'b0;
    end else if(1'b1) begin
      scause_q[31] <= scause_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[30] <= 1'b0;
    end else if(1'b1) begin
      scause_q[30] <= scause_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[29] <= 1'b0;
    end else if(1'b1) begin
      scause_q[29] <= scause_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[28] <= 1'b0;
    end else if(1'b1) begin
      scause_q[28] <= scause_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[27] <= 1'b0;
    end else if(1'b1) begin
      scause_q[27] <= scause_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[26] <= 1'b0;
    end else if(1'b1) begin
      scause_q[26] <= scause_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[25] <= 1'b0;
    end else if(1'b1) begin
      scause_q[25] <= scause_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[24] <= 1'b0;
    end else if(1'b1) begin
      scause_q[24] <= scause_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[23] <= 1'b0;
    end else if(1'b1) begin
      scause_q[23] <= scause_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[22] <= 1'b0;
    end else if(1'b1) begin
      scause_q[22] <= scause_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[21] <= 1'b0;
    end else if(1'b1) begin
      scause_q[21] <= scause_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[20] <= 1'b0;
    end else if(1'b1) begin
      scause_q[20] <= scause_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[19] <= 1'b0;
    end else if(1'b1) begin
      scause_q[19] <= scause_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[18] <= 1'b0;
    end else if(1'b1) begin
      scause_q[18] <= scause_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[17] <= 1'b0;
    end else if(1'b1) begin
      scause_q[17] <= scause_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[16] <= 1'b0;
    end else if(1'b1) begin
      scause_q[16] <= scause_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[15] <= 1'b0;
    end else if(1'b1) begin
      scause_q[15] <= scause_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[14] <= 1'b0;
    end else if(1'b1) begin
      scause_q[14] <= scause_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[13] <= 1'b0;
    end else if(1'b1) begin
      scause_q[13] <= scause_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[12] <= 1'b0;
    end else if(1'b1) begin
      scause_q[12] <= scause_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[11] <= 1'b0;
    end else if(1'b1) begin
      scause_q[11] <= scause_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[10] <= 1'b0;
    end else if(1'b1) begin
      scause_q[10] <= scause_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[9] <= 1'b0;
    end else if(1'b1) begin
      scause_q[9] <= scause_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[8] <= 1'b0;
    end else if(1'b1) begin
      scause_q[8] <= scause_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[7] <= 1'b0;
    end else if(1'b1) begin
      scause_q[7] <= scause_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[6] <= 1'b0;
    end else if(1'b1) begin
      scause_q[6] <= scause_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[5] <= 1'b0;
    end else if(1'b1) begin
      scause_q[5] <= scause_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[4] <= 1'b0;
    end else if(1'b1) begin
      scause_q[4] <= scause_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[3] <= 1'b0;
    end else if(1'b1) begin
      scause_q[3] <= scause_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[2] <= 1'b0;
    end else if(1'b1) begin
      scause_q[2] <= scause_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[1] <= 1'b0;
    end else if(1'b1) begin
      scause_q[1] <= scause_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      scause_q[0] <= 1'b0;
    end else if(1'b1) begin
      scause_q[0] <= scause_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[63] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[63] <= stvec_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[62] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[62] <= stvec_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[61] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[61] <= stvec_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[60] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[60] <= stvec_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[59] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[59] <= stvec_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[58] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[58] <= stvec_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[57] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[57] <= stvec_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[56] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[56] <= stvec_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[55] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[55] <= stvec_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[54] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[54] <= stvec_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[53] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[53] <= stvec_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[52] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[52] <= stvec_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[51] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[51] <= stvec_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[50] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[50] <= stvec_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[49] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[49] <= stvec_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[48] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[48] <= stvec_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[47] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[47] <= stvec_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[46] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[46] <= stvec_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[45] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[45] <= stvec_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[44] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[44] <= stvec_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[43] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[43] <= stvec_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[42] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[42] <= stvec_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[41] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[41] <= stvec_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[40] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[40] <= stvec_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[39] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[39] <= stvec_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[38] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[38] <= stvec_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[37] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[37] <= stvec_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[36] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[36] <= stvec_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[35] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[35] <= stvec_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[34] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[34] <= stvec_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[33] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[33] <= stvec_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[32] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[32] <= stvec_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[31] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[31] <= stvec_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[30] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[30] <= stvec_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[29] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[29] <= stvec_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[28] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[28] <= stvec_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[27] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[27] <= stvec_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[26] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[26] <= stvec_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[25] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[25] <= stvec_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[24] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[24] <= stvec_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[23] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[23] <= stvec_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[22] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[22] <= stvec_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[21] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[21] <= stvec_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[20] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[20] <= stvec_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[19] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[19] <= stvec_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[18] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[18] <= stvec_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[17] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[17] <= stvec_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[16] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[16] <= stvec_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[15] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[15] <= stvec_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[14] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[14] <= stvec_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[13] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[13] <= stvec_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[12] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[12] <= stvec_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[11] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[11] <= stvec_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[10] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[10] <= stvec_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[9] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[9] <= stvec_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[8] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[8] <= stvec_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[7] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[7] <= stvec_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[6] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[6] <= stvec_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[5] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[5] <= stvec_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[4] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[4] <= stvec_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[3] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[3] <= stvec_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[2] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[2] <= stvec_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[1] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[1] <= stvec_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stvec_q[0] <= 1'b0;
    end else if(1'b1) begin
      stvec_q[0] <= stvec_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[63] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[63] <= sscratch_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[62] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[62] <= sscratch_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[61] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[61] <= sscratch_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[60] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[60] <= sscratch_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[59] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[59] <= sscratch_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[58] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[58] <= sscratch_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[57] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[57] <= sscratch_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[56] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[56] <= sscratch_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[55] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[55] <= sscratch_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[54] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[54] <= sscratch_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[53] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[53] <= sscratch_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[52] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[52] <= sscratch_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[51] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[51] <= sscratch_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[50] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[50] <= sscratch_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[49] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[49] <= sscratch_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[48] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[48] <= sscratch_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[47] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[47] <= sscratch_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[46] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[46] <= sscratch_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[45] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[45] <= sscratch_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[44] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[44] <= sscratch_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[43] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[43] <= sscratch_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[42] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[42] <= sscratch_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[41] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[41] <= sscratch_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[40] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[40] <= sscratch_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[39] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[39] <= sscratch_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[38] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[38] <= sscratch_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[37] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[37] <= sscratch_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[36] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[36] <= sscratch_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[35] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[35] <= sscratch_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[34] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[34] <= sscratch_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[33] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[33] <= sscratch_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[32] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[32] <= sscratch_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[31] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[31] <= sscratch_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[30] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[30] <= sscratch_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[29] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[29] <= sscratch_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[28] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[28] <= sscratch_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[27] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[27] <= sscratch_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[26] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[26] <= sscratch_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[25] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[25] <= sscratch_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[24] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[24] <= sscratch_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[23] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[23] <= sscratch_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[22] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[22] <= sscratch_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[21] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[21] <= sscratch_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[20] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[20] <= sscratch_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[19] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[19] <= sscratch_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[18] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[18] <= sscratch_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[17] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[17] <= sscratch_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[16] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[16] <= sscratch_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[15] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[15] <= sscratch_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[14] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[14] <= sscratch_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[13] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[13] <= sscratch_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[12] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[12] <= sscratch_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[11] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[11] <= sscratch_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[10] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[10] <= sscratch_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[9] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[9] <= sscratch_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[8] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[8] <= sscratch_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[7] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[7] <= sscratch_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[6] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[6] <= sscratch_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[5] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[5] <= sscratch_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[4] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[4] <= sscratch_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[3] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[3] <= sscratch_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[2] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[2] <= sscratch_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[1] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[1] <= sscratch_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      sscratch_q[0] <= 1'b0;
    end else if(1'b1) begin
      sscratch_q[0] <= sscratch_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[63] <= 1'b0;
    end else if(1'b1) begin
      stval_q[63] <= stval_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[62] <= 1'b0;
    end else if(1'b1) begin
      stval_q[62] <= stval_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[61] <= 1'b0;
    end else if(1'b1) begin
      stval_q[61] <= stval_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[60] <= 1'b0;
    end else if(1'b1) begin
      stval_q[60] <= stval_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[59] <= 1'b0;
    end else if(1'b1) begin
      stval_q[59] <= stval_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[58] <= 1'b0;
    end else if(1'b1) begin
      stval_q[58] <= stval_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[57] <= 1'b0;
    end else if(1'b1) begin
      stval_q[57] <= stval_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[56] <= 1'b0;
    end else if(1'b1) begin
      stval_q[56] <= stval_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[55] <= 1'b0;
    end else if(1'b1) begin
      stval_q[55] <= stval_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[54] <= 1'b0;
    end else if(1'b1) begin
      stval_q[54] <= stval_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[53] <= 1'b0;
    end else if(1'b1) begin
      stval_q[53] <= stval_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[52] <= 1'b0;
    end else if(1'b1) begin
      stval_q[52] <= stval_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[51] <= 1'b0;
    end else if(1'b1) begin
      stval_q[51] <= stval_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[50] <= 1'b0;
    end else if(1'b1) begin
      stval_q[50] <= stval_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[49] <= 1'b0;
    end else if(1'b1) begin
      stval_q[49] <= stval_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[48] <= 1'b0;
    end else if(1'b1) begin
      stval_q[48] <= stval_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[47] <= 1'b0;
    end else if(1'b1) begin
      stval_q[47] <= stval_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[46] <= 1'b0;
    end else if(1'b1) begin
      stval_q[46] <= stval_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[45] <= 1'b0;
    end else if(1'b1) begin
      stval_q[45] <= stval_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[44] <= 1'b0;
    end else if(1'b1) begin
      stval_q[44] <= stval_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[43] <= 1'b0;
    end else if(1'b1) begin
      stval_q[43] <= stval_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[42] <= 1'b0;
    end else if(1'b1) begin
      stval_q[42] <= stval_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[41] <= 1'b0;
    end else if(1'b1) begin
      stval_q[41] <= stval_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[40] <= 1'b0;
    end else if(1'b1) begin
      stval_q[40] <= stval_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[39] <= 1'b0;
    end else if(1'b1) begin
      stval_q[39] <= stval_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[38] <= 1'b0;
    end else if(1'b1) begin
      stval_q[38] <= stval_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[37] <= 1'b0;
    end else if(1'b1) begin
      stval_q[37] <= stval_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[36] <= 1'b0;
    end else if(1'b1) begin
      stval_q[36] <= stval_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[35] <= 1'b0;
    end else if(1'b1) begin
      stval_q[35] <= stval_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[34] <= 1'b0;
    end else if(1'b1) begin
      stval_q[34] <= stval_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[33] <= 1'b0;
    end else if(1'b1) begin
      stval_q[33] <= stval_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[32] <= 1'b0;
    end else if(1'b1) begin
      stval_q[32] <= stval_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[31] <= 1'b0;
    end else if(1'b1) begin
      stval_q[31] <= stval_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[30] <= 1'b0;
    end else if(1'b1) begin
      stval_q[30] <= stval_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[29] <= 1'b0;
    end else if(1'b1) begin
      stval_q[29] <= stval_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[28] <= 1'b0;
    end else if(1'b1) begin
      stval_q[28] <= stval_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[27] <= 1'b0;
    end else if(1'b1) begin
      stval_q[27] <= stval_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[26] <= 1'b0;
    end else if(1'b1) begin
      stval_q[26] <= stval_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[25] <= 1'b0;
    end else if(1'b1) begin
      stval_q[25] <= stval_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[24] <= 1'b0;
    end else if(1'b1) begin
      stval_q[24] <= stval_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[23] <= 1'b0;
    end else if(1'b1) begin
      stval_q[23] <= stval_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[22] <= 1'b0;
    end else if(1'b1) begin
      stval_q[22] <= stval_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[21] <= 1'b0;
    end else if(1'b1) begin
      stval_q[21] <= stval_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[20] <= 1'b0;
    end else if(1'b1) begin
      stval_q[20] <= stval_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[19] <= 1'b0;
    end else if(1'b1) begin
      stval_q[19] <= stval_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[18] <= 1'b0;
    end else if(1'b1) begin
      stval_q[18] <= stval_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[17] <= 1'b0;
    end else if(1'b1) begin
      stval_q[17] <= stval_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[16] <= 1'b0;
    end else if(1'b1) begin
      stval_q[16] <= stval_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[15] <= 1'b0;
    end else if(1'b1) begin
      stval_q[15] <= stval_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[14] <= 1'b0;
    end else if(1'b1) begin
      stval_q[14] <= stval_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[13] <= 1'b0;
    end else if(1'b1) begin
      stval_q[13] <= stval_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[12] <= 1'b0;
    end else if(1'b1) begin
      stval_q[12] <= stval_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[11] <= 1'b0;
    end else if(1'b1) begin
      stval_q[11] <= stval_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[10] <= 1'b0;
    end else if(1'b1) begin
      stval_q[10] <= stval_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[9] <= 1'b0;
    end else if(1'b1) begin
      stval_q[9] <= stval_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[8] <= 1'b0;
    end else if(1'b1) begin
      stval_q[8] <= stval_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[7] <= 1'b0;
    end else if(1'b1) begin
      stval_q[7] <= stval_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[6] <= 1'b0;
    end else if(1'b1) begin
      stval_q[6] <= stval_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[5] <= 1'b0;
    end else if(1'b1) begin
      stval_q[5] <= stval_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[4] <= 1'b0;
    end else if(1'b1) begin
      stval_q[4] <= stval_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[3] <= 1'b0;
    end else if(1'b1) begin
      stval_q[3] <= stval_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[2] <= 1'b0;
    end else if(1'b1) begin
      stval_q[2] <= stval_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[1] <= 1'b0;
    end else if(1'b1) begin
      stval_q[1] <= stval_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      stval_q[0] <= 1'b0;
    end else if(1'b1) begin
      stval_q[0] <= stval_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_mode__3_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_mode__3_ <= satp_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_mode__2_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_mode__2_ <= satp_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_mode__1_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_mode__1_ <= satp_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_mode__0_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_mode__0_ <= satp_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__15_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__15_ <= satp_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__14_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__14_ <= satp_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__13_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__13_ <= satp_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__12_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__12_ <= satp_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__11_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__11_ <= satp_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__10_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__10_ <= satp_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__9_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__9_ <= satp_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__8_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__8_ <= satp_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__7_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__7_ <= satp_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__6_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__6_ <= satp_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__5_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__5_ <= satp_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__4_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__4_ <= satp_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__3_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__3_ <= satp_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__2_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__2_ <= satp_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_q_asid__1_ <= 1'b0;
    end else if(1'b1) begin
      satp_q_asid__1_ <= satp_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      asid_o[0] <= 1'b0;
    end else if(1'b1) begin
      asid_o[0] <= satp_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[43] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[43] <= satp_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[42] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[42] <= satp_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[41] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[41] <= satp_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[40] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[40] <= satp_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[39] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[39] <= satp_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[38] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[38] <= satp_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[37] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[37] <= satp_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[36] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[36] <= satp_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[35] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[35] <= satp_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[34] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[34] <= satp_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[33] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[33] <= satp_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[32] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[32] <= satp_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[31] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[31] <= satp_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[30] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[30] <= satp_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[29] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[29] <= satp_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[28] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[28] <= satp_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[27] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[27] <= satp_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[26] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[26] <= satp_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[25] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[25] <= satp_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[24] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[24] <= satp_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[23] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[23] <= satp_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[22] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[22] <= satp_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[21] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[21] <= satp_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[20] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[20] <= satp_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[19] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[19] <= satp_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[18] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[18] <= satp_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[17] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[17] <= satp_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[16] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[16] <= satp_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[15] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[15] <= satp_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[14] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[14] <= satp_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[13] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[13] <= satp_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[12] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[12] <= satp_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[11] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[11] <= satp_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[10] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[10] <= satp_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[9] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[9] <= satp_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[8] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[8] <= satp_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[7] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[7] <= satp_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[6] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[6] <= satp_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[5] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[5] <= satp_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[4] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[4] <= satp_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[3] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[3] <= satp_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[2] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[2] <= satp_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[1] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[1] <= satp_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      satp_ppn_o[0] <= 1'b0;
    end else if(1'b1) begin
      satp_ppn_o[0] <= satp_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[63] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[63] <= cycle_d[63];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[62] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[62] <= cycle_d[62];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[61] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[61] <= cycle_d[61];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[60] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[60] <= cycle_d[60];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[59] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[59] <= cycle_d[59];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[58] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[58] <= cycle_d[58];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[57] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[57] <= cycle_d[57];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[56] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[56] <= cycle_d[56];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[55] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[55] <= cycle_d[55];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[54] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[54] <= cycle_d[54];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[53] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[53] <= cycle_d[53];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[52] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[52] <= cycle_d[52];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[51] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[51] <= cycle_d[51];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[50] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[50] <= cycle_d[50];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[49] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[49] <= cycle_d[49];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[48] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[48] <= cycle_d[48];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[47] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[47] <= cycle_d[47];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[46] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[46] <= cycle_d[46];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[45] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[45] <= cycle_d[45];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[44] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[44] <= cycle_d[44];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[43] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[43] <= cycle_d[43];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[42] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[42] <= cycle_d[42];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[41] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[41] <= cycle_d[41];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[40] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[40] <= cycle_d[40];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[39] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[39] <= cycle_d[39];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[38] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[38] <= cycle_d[38];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[37] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[37] <= cycle_d[37];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[36] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[36] <= cycle_d[36];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[35] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[35] <= cycle_d[35];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[34] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[34] <= cycle_d[34];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[33] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[33] <= cycle_d[33];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[32] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[32] <= cycle_d[32];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[31] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[31] <= cycle_d[31];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[30] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[30] <= cycle_d[30];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[29] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[29] <= cycle_d[29];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[28] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[28] <= cycle_d[28];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[27] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[27] <= cycle_d[27];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[26] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[26] <= cycle_d[26];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[25] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[25] <= cycle_d[25];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[24] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[24] <= cycle_d[24];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[23] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[23] <= cycle_d[23];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[22] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[22] <= cycle_d[22];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[21] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[21] <= cycle_d[21];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[20] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[20] <= cycle_d[20];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[19] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[19] <= cycle_d[19];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[18] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[18] <= cycle_d[18];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[17] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[17] <= cycle_d[17];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[16] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[16] <= cycle_d[16];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[15] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[15] <= cycle_d[15];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[14] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[14] <= cycle_d[14];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[13] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[13] <= cycle_d[13];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[12] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[12] <= cycle_d[12];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[11] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[11] <= cycle_d[11];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[10] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[10] <= cycle_d[10];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[9] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[9] <= cycle_d[9];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[8] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[8] <= cycle_d[8];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[7] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[7] <= cycle_d[7];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[6] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[6] <= cycle_d[6];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[5] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[5] <= cycle_d[5];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[4] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[4] <= cycle_d[4];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[3] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[3] <= cycle_d[3];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[2] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[2] <= cycle_d[2];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[1] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[1] <= cycle_d[1];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      cycle_q[0] <= 1'b0;
    end else if(1'b1) begin
      cycle_q[0] <= cycle_d[0];
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[63] <= 1'b0;
    end else if(N5437) begin
      instret_q[63] <= N1292;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[62] <= 1'b0;
    end else if(N5437) begin
      instret_q[62] <= N1291;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[61] <= 1'b0;
    end else if(N5437) begin
      instret_q[61] <= N1290;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[60] <= 1'b0;
    end else if(N5437) begin
      instret_q[60] <= N1289;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[59] <= 1'b0;
    end else if(N5437) begin
      instret_q[59] <= N1288;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[58] <= 1'b0;
    end else if(N5437) begin
      instret_q[58] <= N1287;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[57] <= 1'b0;
    end else if(N5437) begin
      instret_q[57] <= N1286;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[56] <= 1'b0;
    end else if(N5437) begin
      instret_q[56] <= N1285;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[55] <= 1'b0;
    end else if(N5437) begin
      instret_q[55] <= N1284;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[54] <= 1'b0;
    end else if(N5437) begin
      instret_q[54] <= N1283;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[53] <= 1'b0;
    end else if(N5437) begin
      instret_q[53] <= N1282;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[52] <= 1'b0;
    end else if(N5437) begin
      instret_q[52] <= N1281;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[51] <= 1'b0;
    end else if(N5437) begin
      instret_q[51] <= N1280;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[50] <= 1'b0;
    end else if(N5437) begin
      instret_q[50] <= N1279;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[49] <= 1'b0;
    end else if(N5437) begin
      instret_q[49] <= N1278;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[48] <= 1'b0;
    end else if(N5437) begin
      instret_q[48] <= N1277;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[47] <= 1'b0;
    end else if(N5437) begin
      instret_q[47] <= N1276;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[46] <= 1'b0;
    end else if(N5437) begin
      instret_q[46] <= N1275;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[45] <= 1'b0;
    end else if(N5437) begin
      instret_q[45] <= N1274;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[44] <= 1'b0;
    end else if(N5437) begin
      instret_q[44] <= N1273;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[43] <= 1'b0;
    end else if(N5437) begin
      instret_q[43] <= N1272;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[42] <= 1'b0;
    end else if(N5437) begin
      instret_q[42] <= N1271;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[41] <= 1'b0;
    end else if(N5437) begin
      instret_q[41] <= N1270;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[40] <= 1'b0;
    end else if(N5437) begin
      instret_q[40] <= N1269;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[39] <= 1'b0;
    end else if(N5437) begin
      instret_q[39] <= N1268;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[38] <= 1'b0;
    end else if(N5437) begin
      instret_q[38] <= N1267;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[37] <= 1'b0;
    end else if(N5437) begin
      instret_q[37] <= N1266;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[36] <= 1'b0;
    end else if(N5437) begin
      instret_q[36] <= N1265;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[35] <= 1'b0;
    end else if(N5437) begin
      instret_q[35] <= N1264;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[34] <= 1'b0;
    end else if(N5437) begin
      instret_q[34] <= N1263;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[33] <= 1'b0;
    end else if(N5437) begin
      instret_q[33] <= N1262;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[32] <= 1'b0;
    end else if(N5437) begin
      instret_q[32] <= N1261;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[31] <= 1'b0;
    end else if(N5437) begin
      instret_q[31] <= N1260;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[30] <= 1'b0;
    end else if(N5437) begin
      instret_q[30] <= N1259;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[29] <= 1'b0;
    end else if(N5437) begin
      instret_q[29] <= N1258;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[28] <= 1'b0;
    end else if(N5437) begin
      instret_q[28] <= N1257;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[27] <= 1'b0;
    end else if(N5437) begin
      instret_q[27] <= N1256;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[26] <= 1'b0;
    end else if(N5437) begin
      instret_q[26] <= N1255;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[25] <= 1'b0;
    end else if(N5437) begin
      instret_q[25] <= N1254;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[24] <= 1'b0;
    end else if(N5437) begin
      instret_q[24] <= N1253;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[23] <= 1'b0;
    end else if(N5437) begin
      instret_q[23] <= N1252;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[22] <= 1'b0;
    end else if(N5437) begin
      instret_q[22] <= N1251;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[21] <= 1'b0;
    end else if(N5437) begin
      instret_q[21] <= N1250;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[20] <= 1'b0;
    end else if(N5437) begin
      instret_q[20] <= N1249;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[19] <= 1'b0;
    end else if(N5437) begin
      instret_q[19] <= N1248;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[18] <= 1'b0;
    end else if(N5437) begin
      instret_q[18] <= N1247;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[17] <= 1'b0;
    end else if(N5437) begin
      instret_q[17] <= N1246;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[16] <= 1'b0;
    end else if(N5437) begin
      instret_q[16] <= N1245;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[15] <= 1'b0;
    end else if(N5437) begin
      instret_q[15] <= N1244;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[14] <= 1'b0;
    end else if(N5437) begin
      instret_q[14] <= N1243;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[13] <= 1'b0;
    end else if(N5437) begin
      instret_q[13] <= N1242;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[12] <= 1'b0;
    end else if(N5437) begin
      instret_q[12] <= N1241;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[11] <= 1'b0;
    end else if(N5437) begin
      instret_q[11] <= N1240;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[10] <= 1'b0;
    end else if(N5437) begin
      instret_q[10] <= N1239;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[9] <= 1'b0;
    end else if(N5437) begin
      instret_q[9] <= N1238;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[8] <= 1'b0;
    end else if(N5437) begin
      instret_q[8] <= N1237;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[7] <= 1'b0;
    end else if(N5437) begin
      instret_q[7] <= N1236;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[6] <= 1'b0;
    end else if(N5437) begin
      instret_q[6] <= N1235;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[5] <= 1'b0;
    end else if(N5437) begin
      instret_q[5] <= N1234;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[4] <= 1'b0;
    end else if(N5437) begin
      instret_q[4] <= N1233;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[3] <= 1'b0;
    end else if(N5437) begin
      instret_q[3] <= N1232;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[2] <= 1'b0;
    end else if(N5437) begin
      instret_q[2] <= N1231;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[1] <= 1'b0;
    end else if(N5437) begin
      instret_q[1] <= N1230;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      instret_q[0] <= 1'b0;
    end else if(N5437) begin
      instret_q[0] <= N1229;
    end 
  end


  always @(posedge clk_i or posedge N5436) begin
    if(N5436) begin
      en_ld_st_translation_o <= 1'b0;
    end else if(1'b1) begin
      en_ld_st_translation_o <= en_ld_st_translation_d;
    end 
  end

  assign N5438 = ~ex_i[66];
  assign N5439 = ~ex_i[65];
  assign N5440 = ex_i[127] | ex_i[128];
  assign N5441 = ex_i[126] | N5440;
  assign N5442 = ex_i[125] | N5441;
  assign N5443 = ex_i[124] | N5442;
  assign N5444 = ex_i[123] | N5443;
  assign N5445 = ex_i[122] | N5444;
  assign N5446 = ex_i[121] | N5445;
  assign N5447 = ex_i[120] | N5446;
  assign N5448 = ex_i[119] | N5447;
  assign N5449 = ex_i[118] | N5448;
  assign N5450 = ex_i[117] | N5449;
  assign N5451 = ex_i[116] | N5450;
  assign N5452 = ex_i[115] | N5451;
  assign N5453 = ex_i[114] | N5452;
  assign N5454 = ex_i[113] | N5453;
  assign N5455 = ex_i[112] | N5454;
  assign N5456 = ex_i[111] | N5455;
  assign N5457 = ex_i[110] | N5456;
  assign N5458 = ex_i[109] | N5457;
  assign N5459 = ex_i[108] | N5458;
  assign N5460 = ex_i[107] | N5459;
  assign N5461 = ex_i[106] | N5460;
  assign N5462 = ex_i[105] | N5461;
  assign N5463 = ex_i[104] | N5462;
  assign N5464 = ex_i[103] | N5463;
  assign N5465 = ex_i[102] | N5464;
  assign N5466 = ex_i[101] | N5465;
  assign N5467 = ex_i[100] | N5466;
  assign N5468 = ex_i[99] | N5467;
  assign N5469 = ex_i[98] | N5468;
  assign N5470 = ex_i[97] | N5469;
  assign N5471 = ex_i[96] | N5470;
  assign N5472 = ex_i[95] | N5471;
  assign N5473 = ex_i[94] | N5472;
  assign N5474 = ex_i[93] | N5473;
  assign N5475 = ex_i[92] | N5474;
  assign N5476 = ex_i[91] | N5475;
  assign N5477 = ex_i[90] | N5476;
  assign N5478 = ex_i[89] | N5477;
  assign N5479 = ex_i[88] | N5478;
  assign N5480 = ex_i[87] | N5479;
  assign N5481 = ex_i[86] | N5480;
  assign N5482 = ex_i[85] | N5481;
  assign N5483 = ex_i[84] | N5482;
  assign N5484 = ex_i[83] | N5483;
  assign N5485 = ex_i[82] | N5484;
  assign N5486 = ex_i[81] | N5485;
  assign N5487 = ex_i[80] | N5486;
  assign N5488 = ex_i[79] | N5487;
  assign N5489 = ex_i[78] | N5488;
  assign N5490 = ex_i[77] | N5489;
  assign N5491 = ex_i[76] | N5490;
  assign N5492 = ex_i[75] | N5491;
  assign N5493 = ex_i[74] | N5492;
  assign N5494 = ex_i[73] | N5493;
  assign N5495 = ex_i[72] | N5494;
  assign N5496 = ex_i[71] | N5495;
  assign N5497 = ex_i[70] | N5496;
  assign N5498 = ex_i[69] | N5497;
  assign N5499 = ex_i[68] | N5498;
  assign N5500 = ex_i[67] | N5499;
  assign N5501 = N5438 | N5500;
  assign N5502 = N5439 | N5501;
  assign N5503 = ~N5502;
  assign N5504 = ~satp_q_mode__3_;
  assign N5505 = satp_q_mode__2_ | N5504;
  assign N5506 = satp_q_mode__1_ | N5505;
  assign N5507 = satp_q_mode__0_ | N5506;
  assign N5508 = ~N5507;
  assign N5509 = mstatus_q_mpp__0_ & mstatus_q_mpp__1_;
  assign N5510 = ~N5509;
  assign N5511 = ~csr_op_i[4];
  assign N5512 = ~csr_op_i[3];
  assign N5513 = ~csr_op_i[1];
  assign N5514 = csr_op_i[5] | csr_op_i[6];
  assign N5515 = N5511 | N5514;
  assign N5516 = N5512 | N5515;
  assign N5517 = csr_op_i[2] | N5516;
  assign N5518 = N5513 | N5517;
  assign N5519 = csr_op_i[0] | N5518;
  assign N5520 = ~N5519;
  assign N5521 = ~N4160;
  assign N5522 = satp_q_mode__2_ | N5504;
  assign N5523 = satp_q_mode__1_ | N5522;
  assign N5524 = satp_q_mode__0_ | N5523;
  assign N5525 = ~N5524;
  assign N5526 = priv_lvl_o[0] & priv_lvl_o[1];
  assign N5527 = ~N5526;
  assign N5528 = csr_wdata[62] | csr_wdata[63];
  assign N5529 = csr_wdata[61] | N5528;
  assign N5530 = csr_wdata[60] | N5529;
  assign N5531 = ~N5530;
  assign N5532 = ~csr_wdata[63];
  assign N5533 = csr_wdata[62] | N5532;
  assign N5534 = csr_wdata[61] | N5533;
  assign N5535 = csr_wdata[60] | N5534;
  assign N5536 = ~N5535;
  assign N5537 = ~trap_to_priv_lvl[1];
  assign N5538 = ~commit_instr_i[293];
  assign N5539 = N5538 | commit_instr_i[294];
  assign N5540 = commit_instr_i[292] | N5539;
  assign N5541 = commit_instr_i[291] | N5540;
  assign N5542 = ~N5541;
  assign N5543 = ~priv_lvl_o[0];
  assign N5544 = N5543 | priv_lvl_o[1];
  assign N5545 = ~N5544;
  assign N5546 = priv_lvl_o[0] | priv_lvl_o[1];
  assign N5547 = ~N5546;
  assign N5548 = ~csr_addr_i[10];
  assign N5549 = ~csr_addr_i[9];
  assign N5550 = ~csr_addr_i[8];
  assign N5551 = ~csr_addr_i[7];
  assign N5552 = ~csr_addr_i[5];
  assign N5553 = ~csr_addr_i[4];
  assign N5554 = N5548 | csr_addr_i[11];
  assign N5555 = N5549 | N5554;
  assign N5556 = N5550 | N5555;
  assign N5557 = N5551 | N5556;
  assign N5558 = csr_addr_i[6] | N5557;
  assign N5559 = N5552 | N5558;
  assign N5560 = N5553 | N5559;
  assign N5561 = ~N5560;
  assign N5562 = priv_lvl_o[0] & priv_lvl_o[1];
  assign N5563 = priv_lvl_o[0] & priv_lvl_o[1];
  assign N5564 = priv_lvl_o[0] & priv_lvl_o[1];
  assign N5565 = ~N5564;
  assign N5566 = fs_o[0] | fs_o[1];
  assign N5567 = ~N5566;
  assign N5568 = fs_o[0] | fs_o[1];
  assign N5569 = ~N5568;
  assign N5570 = fs_o[0] | fs_o[1];
  assign N5571 = ~N5570;
  assign N5572 = fs_o[0] | fs_o[1];
  assign N5573 = ~N5572;
  assign N5574 = fs_o[0] | fs_o[1];
  assign N5575 = ~N5574;
  assign N5576 = fs_o[0] | fs_o[1];
  assign N5577 = ~N5576;
  assign N5578 = fs_o[0] | fs_o[1];
  assign N5579 = ~N5578;
  assign N5580 = fs_o[0] | fs_o[1];
  assign N5581 = ~N5580;
  assign N5582 = N5543 | priv_lvl_o[1];
  assign N5583 = ~N5582;
  assign N5584 = N5543 | priv_lvl_o[1];
  assign N5585 = ~N5584;
  assign { N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422 } = boot_addr_i + { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293 } = cycle_q + 1'b1;
  assign { N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035 } = instret_q + 1'b1;
  assign { N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719 } = commit_instr_i[361:298] + { N4718, commit_instr_i[0:0], 1'b0 };
  assign { N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165 } = { N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099 } + 1'b1;
  assign { N751, N750, N749, N748, N747 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N2)? fflags_o : 1'b0;
  assign N1 = N5575;
  assign N2 = N5574;
  assign { N754, N753, N752 } = (N3)? { 1'b0, 1'b0, 1'b0 } : 
                                (N4)? frm_o : 1'b0;
  assign N3 = N5577;
  assign N4 = N5576;
  assign { N762, N761, N760, N759, N758, N757, N756, N755 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                              (N6)? { frm_o, fflags_o } : 1'b0;
  assign N5 = N5579;
  assign N6 = N5578;
  assign { N769, N768, N767, N766, N765, N764, N763 } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N8)? fprec_o : 1'b0;
  assign N7 = N5581;
  assign N8 = N5580;
  assign { N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900 } = (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N899)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 1'b0;
  assign N9 = N898;
  assign { N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N751, N750, N749, N748, N747 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N754, N753, N752 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N762, N761, N760, N759, N758, N757, N756, N755 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N769, N768, N767, N766, N765, N764, N763 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N15)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N16)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N17)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N22)? { mstatus_q_sd_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mstatus_q_uxl__1_, mstatus_q_uxl__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mxr_o, sum_o, 1'b0, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, 1'b0, 1'b0, 1'b0, 1'b0, mstatus_q_spp_, 1'b0, 1'b0, mstatus_q_spie_, mstatus_q_upie_, 1'b0, 1'b0, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N23)? { N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N24)? { N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N25)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N27)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N28)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N29)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N30)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N31)? { N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N32)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_sxl__1_, mstatus_q_sxl__0_, mstatus_q_uxl__1_, mstatus_q_uxl__0_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N33)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N34)? { medeleg_d[63:16], medeleg_q_15, medeleg_d[14:14], medeleg_q, medeleg_d[11:9], medeleg_q_8, medeleg_d[7:4], medeleg_q_3, medeleg_d[2:1], medeleg_q_0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N35)? { mideleg_d[63:10], mideleg_q[9:9], mideleg_d[8:6], mideleg_q_5, mideleg_d[4:2], mideleg_q_1, mideleg_d[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N36)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N37)? mtvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N39)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N40)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N41)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N42)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N43)? { mip_d, mip_q[11:11], mip_d_10, mip_q_9, mip_d_8, mip_q_7, mip_d_6, mip_q_5, mip_d_4, mip_q_3, mip_d_2, mip_q_1, mip_d_0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N44)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N45)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N47)? hart_id_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N48)? cycle_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N49)? instret_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N50)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N51)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N52)? cycle_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N53)? instret_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N54)? perf_data_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                          (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N179;
  assign N11 = N188;
  assign N12 = N196;
  assign N13 = N206;
  assign N14 = N215;
  assign N15 = N223;
  assign N16 = N231;
  assign N17 = N239;
  assign N18 = N247;
  assign N19 = N255;
  assign N20 = N263;
  assign N21 = N271;
  assign N22 = N279;
  assign N23 = N288;
  assign N24 = N296;
  assign N25 = N304;
  assign N26 = N312;
  assign N27 = N320;
  assign N28 = N328;
  assign N29 = N336;
  assign N30 = N344;
  assign N31 = N352;
  assign N32 = N360;
  assign N33 = N368;
  assign N34 = N376;
  assign N35 = N384;
  assign N36 = N392;
  assign N37 = N400;
  assign N38 = N408;
  assign N39 = N416;
  assign N40 = N424;
  assign N41 = N432;
  assign N42 = N440;
  assign N43 = N448;
  assign N44 = N457;
  assign N45 = N465;
  assign N46 = N473;
  assign N47 = N481;
  assign N48 = N490;
  assign N49 = N498;
  assign N50 = N506;
  assign N51 = N514;
  assign N52 = N522;
  assign N53 = N530;
  assign N54 = N630;
  assign N55 = N746;
  assign N1028 = (N10)? N5575 : 
                 (N11)? N5577 : 
                 (N12)? N5579 : 
                 (N13)? N5581 : 
                 (N14)? 1'b0 : 
                 (N15)? 1'b0 : 
                 (N16)? 1'b0 : 
                 (N17)? 1'b0 : 
                 (N18)? 1'b0 : 
                 (N19)? 1'b0 : 
                 (N20)? 1'b0 : 
                 (N21)? 1'b0 : 
                 (N22)? 1'b0 : 
                 (N23)? 1'b0 : 
                 (N24)? 1'b0 : 
                 (N25)? 1'b0 : 
                 (N26)? 1'b0 : 
                 (N27)? 1'b0 : 
                 (N28)? 1'b0 : 
                 (N29)? 1'b0 : 
                 (N30)? 1'b0 : 
                 (N31)? N898 : 
                 (N32)? 1'b0 : 
                 (N33)? 1'b0 : 
                 (N34)? 1'b0 : 
                 (N35)? 1'b0 : 
                 (N36)? 1'b0 : 
                 (N37)? 1'b0 : 
                 (N38)? 1'b0 : 
                 (N39)? 1'b0 : 
                 (N40)? 1'b0 : 
                 (N41)? 1'b0 : 
                 (N42)? 1'b0 : 
                 (N43)? 1'b0 : 
                 (N44)? 1'b0 : 
                 (N45)? 1'b0 : 
                 (N46)? 1'b0 : 
                 (N47)? 1'b0 : 
                 (N48)? 1'b0 : 
                 (N49)? 1'b0 : 
                 (N50)? 1'b0 : 
                 (N51)? 1'b0 : 
                 (N52)? 1'b0 : 
                 (N53)? 1'b0 : 
                 (N54)? 1'b0 : 
                 (N55)? 1'b1 : 1'b0;
  assign { csr_rdata_o[63:10], csr_rdata[9:9], csr_rdata_o[8:0] } = (N56)? { N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964 } : 
                                                                    (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = csr_read;
  assign N57 = N169;
  assign read_access_exception = (N56)? N1028 : 
                                 (N57)? 1'b0 : 1'b0;
  assign { N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099 } = (N58)? { N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1034)? instret_q : 1'b0;
  assign N58 = N1033;
  assign { N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229 } = (N59)? { N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1164)? { N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099 } : 1'b0;
  assign N59 = N1163;
  assign { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } = (N60)? { N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N61)? cycle_q : 1'b0;
  assign N60 = N1030;
  assign N61 = debug_mode_o;
  assign { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } = (N62)? { N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N63)? mtvec_q : 1'b0;
  assign N62 = mtvec_rst_load_q;
  assign N63 = N1421;
  assign { N1990, N1989, N1988, N1987, N1986 } = (N64)? fflags_o : 
                                                 (N65)? csr_wdata[4:0] : 1'b0;
  assign N64 = N5567;
  assign N65 = N5566;
  assign { N1993, N1992, N1991 } = (N66)? frm_o : 
                                   (N67)? csr_wdata[2:0] : 1'b0;
  assign N66 = N5569;
  assign N67 = N5568;
  assign { N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994 } = (N68)? { frm_o, fflags_o } : 
                                                                      (N69)? csr_wdata[7:0] : 1'b0;
  assign N68 = N5571;
  assign N69 = N5570;
  assign { N2008, N2007, N2006, N2005, N2004, N2003, N2002 } = (N70)? fprec_o : 
                                                               (N71)? csr_wdata[6:0] : 1'b0;
  assign N70 = N5573;
  assign N71 = N5572;
  assign { N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078 } = (N72)? { csr_wdata[63:60], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, csr_wdata[44:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2077)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 1'b0;
  assign N72 = N2076;
  assign { N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142 } = (N73)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2075)? { N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078 } : 1'b0;
  assign N73 = N2074;
  assign { N2212, N2211, N2210, N2209, N2208, N2207 } = (N74)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2206)? csr_wdata[7:2] : 1'b0;
  assign N74 = csr_wdata[0];
  assign N2213 = (N75)? N5566 : 
                 (N76)? N5568 : 
                 (N77)? N5570 : 
                 (N78)? N5572 : 
                 (N79)? 1'b0 : 
                 (N80)? 1'b0 : 
                 (N81)? 1'b0 : 
                 (N82)? 1'b0 : 
                 (N83)? 1'b0 : 
                 (N84)? 1'b0 : 
                 (N85)? 1'b0 : 
                 (N86)? 1'b0 : 
                 (N87)? 1'b1 : 
                 (N88)? 1'b0 : 
                 (N89)? 1'b0 : 
                 (N90)? 1'b0 : 
                 (N91)? 1'b0 : 
                 (N92)? 1'b0 : 
                 (N93)? 1'b0 : 
                 (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b1 : 
                 (N97)? 1'b1 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N102)? 1'b0 : 
                 (N103)? 1'b0 : 
                 (N104)? 1'b0 : 
                 (N105)? 1'b0 : 
                 (N106)? 1'b0 : 
                 (N107)? 1'b0 : 
                 (N108)? 1'b0 : 
                 (N109)? 1'b0 : 
                 (N110)? 1'b0 : 
                 (N111)? 1'b0 : 
                 (N112)? 1'b0 : 
                 (N113)? 1'b0 : 
                 (N1985)? 1'b0 : 1'b0;
  assign N75 = N1558;
  assign N76 = N1566;
  assign N77 = N1574;
  assign N78 = N1582;
  assign N79 = N1590;
  assign N80 = N1598;
  assign N81 = N1606;
  assign N82 = N1614;
  assign N83 = N1622;
  assign N84 = N1630;
  assign N85 = N1638;
  assign N86 = N1646;
  assign N87 = N1654;
  assign N88 = N1662;
  assign N89 = N1670;
  assign N90 = N1678;
  assign N91 = N1686;
  assign N92 = N1694;
  assign N93 = N1702;
  assign N94 = N1710;
  assign N95 = N1718;
  assign N96 = N1726;
  assign N97 = N1734;
  assign N98 = N1742;
  assign N99 = N1750;
  assign N100 = N1758;
  assign N101 = N1766;
  assign N102 = N1774;
  assign N103 = N1782;
  assign N104 = N1790;
  assign N105 = N1798;
  assign N106 = N1806;
  assign N107 = N1814;
  assign N108 = N1822;
  assign N109 = N1830;
  assign N110 = N1838;
  assign N111 = N1846;
  assign N112 = N1856;
  assign N113 = N1946;
  assign N2214 = (N75)? N5567 : 
                 (N76)? N5569 : 
                 (N77)? N5571 : 
                 (N78)? N5573 : 
                 (N79)? 1'b0 : 
                 (N80)? 1'b0 : 
                 (N81)? 1'b0 : 
                 (N82)? 1'b0 : 
                 (N83)? 1'b0 : 
                 (N84)? 1'b0 : 
                 (N85)? 1'b0 : 
                 (N86)? 1'b0 : 
                 (N87)? 1'b0 : 
                 (N88)? 1'b0 : 
                 (N89)? 1'b0 : 
                 (N90)? 1'b0 : 
                 (N91)? 1'b0 : 
                 (N92)? 1'b0 : 
                 (N93)? 1'b0 : 
                 (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? N2074 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N102)? 1'b0 : 
                 (N103)? 1'b0 : 
                 (N104)? 1'b0 : 
                 (N105)? 1'b0 : 
                 (N106)? 1'b0 : 
                 (N107)? 1'b0 : 
                 (N108)? 1'b0 : 
                 (N109)? 1'b0 : 
                 (N110)? 1'b0 : 
                 (N111)? 1'b0 : 
                 (N112)? 1'b0 : 
                 (N113)? 1'b0 : 
                 (N1985)? 1'b1 : 1'b0;
  assign { N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215 } = (N75)? { frm_o, N1990, N1989, N1988, N1987, N1986 } : 
                                                                      (N76)? { N1993, N1992, N1991, fflags_o } : 
                                                                      (N77)? { N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994 } : 
                                                                      (N78)? { frm_o, fflags_o } : 
                                                                      (N79)? { frm_o, fflags_o } : 
                                                                      (N80)? { frm_o, fflags_o } : 
                                                                      (N81)? { frm_o, fflags_o } : 
                                                                      (N82)? { frm_o, fflags_o } : 
                                                                      (N83)? { frm_o, fflags_o } : 
                                                                      (N84)? { frm_o, fflags_o } : 
                                                                      (N85)? { frm_o, fflags_o } : 
                                                                      (N86)? { frm_o, fflags_o } : 
                                                                      (N87)? { frm_o, fflags_o } : 
                                                                      (N88)? { frm_o, fflags_o } : 
                                                                      (N89)? { frm_o, fflags_o } : 
                                                                      (N90)? { frm_o, fflags_o } : 
                                                                      (N91)? { frm_o, fflags_o } : 
                                                                      (N92)? { frm_o, fflags_o } : 
                                                                      (N93)? { frm_o, fflags_o } : 
                                                                      (N94)? { frm_o, fflags_o } : 
                                                                      (N95)? { frm_o, fflags_o } : 
                                                                      (N96)? { frm_o, fflags_o } : 
                                                                      (N97)? { frm_o, fflags_o } : 
                                                                      (N98)? { frm_o, fflags_o } : 
                                                                      (N99)? { frm_o, fflags_o } : 
                                                                      (N100)? { frm_o, fflags_o } : 
                                                                      (N101)? { frm_o, fflags_o } : 
                                                                      (N102)? { frm_o, fflags_o } : 
                                                                      (N103)? { frm_o, fflags_o } : 
                                                                      (N104)? { frm_o, fflags_o } : 
                                                                      (N105)? { frm_o, fflags_o } : 
                                                                      (N106)? { frm_o, fflags_o } : 
                                                                      (N107)? { frm_o, fflags_o } : 
                                                                      (N108)? { frm_o, fflags_o } : 
                                                                      (N109)? { frm_o, fflags_o } : 
                                                                      (N110)? { frm_o, fflags_o } : 
                                                                      (N111)? { frm_o, fflags_o } : 
                                                                      (N112)? { frm_o, fflags_o } : 
                                                                      (N113)? { frm_o, fflags_o } : 
                                                                      (N1985)? { frm_o, fflags_o } : 1'b0;
  assign { N2230, N2229, N2228, N2227, N2226, N2225, N2224 } = (N78)? { N2008, N2007, N2006, N2005, N2004, N2003, N2002 } : 
                                                               (N2223)? fprec_o : 1'b0;
  assign { N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231 } = (N75)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N76)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N77)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N78)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N79)? { 1'b0, 1'b1, 1'b0, 1'b0, csr_wdata[27:11], 1'b0, 1'b0, csr_wdata[8:4], 1'b0, csr_wdata[2:2], priv_lvl_q } : 
                                                                                                                                                                                                                                              (N80)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N81)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N82)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N83)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N84)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N85)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N86)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N87)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N88)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N89)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N90)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N91)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N92)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N93)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N94)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N95)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N96)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N97)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N98)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N99)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N100)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N101)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N102)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N103)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N104)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N105)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N106)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N107)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N108)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N109)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N110)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N111)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N112)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N113)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                                                              (N1985)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 1'b0;
  assign { N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263 } = (N75)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? dpc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? dpc_q : 1'b0;
  assign { N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327 } = (N75)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? dscratch0_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? dscratch0_q : 1'b0;
  assign { N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391 } = (N75)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? dscratch1_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? dscratch1_q : 1'b0;
  assign { N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455 } = (N75)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N76)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N77)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N78)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N79)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N80)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N81)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N82)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N83)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N84)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N85)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N86)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N87)? { N1031, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, csr_wdata[19:18], mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, 1'b0, 1'b0, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, csr_wdata[8:8], mstatus_q_mpie_, mstatus_q_wpri1_, csr_wdata[5:5], mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, csr_wdata[1:1], mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N88)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N89)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N90)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N91)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N92)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N93)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N94)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N95)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N96)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N97)? { N1031, csr_wdata[62:36], csr_wdata[31:17], 1'b0, 1'b0, 1'b0, 1'b0, csr_wdata[12:5], 1'b0, csr_wdata[3:1], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N98)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N99)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N100)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N101)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N102)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N103)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N104)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N105)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N106)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N107)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N108)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N109)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N110)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N111)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N112)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N113)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N1985)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 1'b0;
  assign { N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515 } = (N75)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { mie_q[63:10], csr_wdata[9:9], mie_q[8:8], csr_wdata[7:7], mie_q[6:6], csr_wdata[5:5], mie_q[4:4], csr_wdata[3:3], mie_q[2:2], csr_wdata[1:1], mie_q[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? mie_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? mie_q : 1'b0;
  assign { N2581, N2580, N2579 } = (N75)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N76)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N77)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N78)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N79)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N80)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N81)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N82)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N83)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N84)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N85)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N86)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N87)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N88)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N89)? { mip_q_9, mip_q_5, N2073 } : 
                                   (N90)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N91)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N92)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N93)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N94)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N95)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N96)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N97)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N98)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N99)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N100)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N101)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N102)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N103)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N104)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N105)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N106)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N107)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N108)? { csr_wdata[9:9], csr_wdata[5:5], csr_wdata[1:1] } : 
                                   (N109)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N110)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N111)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N112)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N113)? { mip_q_9, mip_q_5, mip_q_1 } : 
                                   (N1985)? { mip_q_9, mip_q_5, mip_q_1 } : 1'b0;
  assign { N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582 } = (N75)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { csr_wdata[63:2], 1'b0, csr_wdata[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? stvec_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? stvec_q : 1'b0;
  assign { N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646 } = (N75)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? sscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? sscratch_q : 1'b0;
  assign { N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710 } = (N75)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { csr_wdata[63:1], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? sepc_q : 1'b0;
  assign { N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774 } = (N75)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? scause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? scause_q : 1'b0;
  assign { N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838 } = (N75)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? stval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? stval_q : 1'b0;
  assign { N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902 } = (N75)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 1'b0;
  assign { N2971, N2970, N2969, N2968, N2967, N2966 } = (N75)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N76)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N77)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N78)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N79)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N80)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N81)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N82)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N83)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N84)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N85)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N86)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N87)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N88)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N89)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N90)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N91)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N92)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N93)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N94)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N95)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N96)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N97)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N98)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N99)? { csr_wdata[15:15], csr_wdata[13:12], csr_wdata[8:8], csr_wdata[3:3], csr_wdata[0:0] } : 
                                                        (N100)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N101)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N102)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N103)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N104)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N105)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N106)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N107)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N108)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N109)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N110)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N111)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N112)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N113)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 
                                                        (N1985)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 1'b0;
  assign { N2974, N2973, N2972 } = (N75)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N76)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N77)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N78)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N79)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N80)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N81)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N82)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N83)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N84)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N85)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N86)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N87)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N88)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N89)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N90)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N91)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N92)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N93)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N94)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N95)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N96)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N97)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N98)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N99)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N100)? { csr_wdata[9:9], csr_wdata[5:5], csr_wdata[1:1] } : 
                                   (N101)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N102)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N103)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N104)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N105)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N106)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N107)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N108)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N109)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N110)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N111)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N112)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N113)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 
                                   (N1985)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 1'b0;
  assign { N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975 } = (N75)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { csr_wdata[63:8], N2212, N2211, N2210, N2209, N2208, N2207, 1'b0, csr_wdata[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 1'b0;
  assign { N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039 } = (N75)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? mscratch_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? mscratch_q : 1'b0;
  assign { N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103 } = (N75)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { csr_wdata[63:1], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? mepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? mepc_q : 1'b0;
  assign { N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167 } = (N75)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? mcause_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? mcause_q : 1'b0;
  assign { N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231 } = (N75)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? mtval_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? mtval_q : 1'b0;
  assign { N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295 } = (N75)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 1'b0;
  assign { N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359 } = (N75)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, csr_wdata[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? { dcache_q, dcache_en_o } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? { dcache_q, dcache_en_o } : 1'b0;
  assign { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423 } = (N75)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, csr_wdata[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? icache_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? icache_q : 1'b0;
  assign { N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487 } = (N75)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N77)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N79)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N80)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N81)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N83)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N85)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N87)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N92)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N93)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N95)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N97)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N98)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N99)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N101)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N103)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N104)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N107)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N109)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N110)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N113)? csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1985)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3551 = (N75)? 1'b0 : 
                 (N76)? 1'b0 : 
                 (N77)? 1'b0 : 
                 (N78)? 1'b0 : 
                 (N79)? 1'b0 : 
                 (N80)? 1'b0 : 
                 (N81)? 1'b0 : 
                 (N82)? 1'b0 : 
                 (N83)? 1'b0 : 
                 (N84)? 1'b0 : 
                 (N85)? 1'b0 : 
                 (N86)? 1'b0 : 
                 (N87)? 1'b0 : 
                 (N88)? 1'b0 : 
                 (N89)? 1'b0 : 
                 (N90)? 1'b0 : 
                 (N91)? 1'b0 : 
                 (N92)? 1'b0 : 
                 (N93)? 1'b0 : 
                 (N94)? 1'b0 : 
                 (N95)? 1'b0 : 
                 (N96)? 1'b0 : 
                 (N97)? 1'b0 : 
                 (N98)? 1'b0 : 
                 (N99)? 1'b0 : 
                 (N100)? 1'b0 : 
                 (N101)? 1'b0 : 
                 (N102)? 1'b0 : 
                 (N103)? 1'b0 : 
                 (N104)? 1'b0 : 
                 (N105)? 1'b0 : 
                 (N106)? 1'b0 : 
                 (N107)? 1'b0 : 
                 (N108)? 1'b0 : 
                 (N109)? 1'b0 : 
                 (N110)? 1'b0 : 
                 (N111)? 1'b0 : 
                 (N112)? 1'b0 : 
                 (N113)? 1'b1 : 
                 (N1985)? 1'b0 : 1'b0;
  assign perf_data_o = (N114)? { N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487 } : 
                       (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N114 = csr_we;
  assign N115 = N1550;
  assign perf_we_o = (N114)? N3551 : 
                     (N115)? 1'b0 : 1'b0;
  assign N3552 = (N114)? N2213 : 
                 (N115)? 1'b0 : 1'b0;
  assign update_access_exception = (N114)? N2214 : 
                                   (N115)? 1'b0 : 1'b0;
  assign { fcsr_d_fprec__6_, fcsr_d_fprec__5_, fcsr_d_fprec__4_, fcsr_d_fprec__3_, fcsr_d_fprec__2_, fcsr_d_fprec__1_, fcsr_d_fprec__0_, fcsr_d_frm__2_, fcsr_d_frm__1_, fcsr_d_frm__0_, N3557, N3556, N3555, N3554, N3553 } = (N114)? { N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215 } : 
                                                                                                                                                                                                                               (N115)? { fprec_o, frm_o, fflags_o } : 1'b0;
  assign { dcsr_d[31:9], N3562, N3561, N3560, dcsr_d[5:2], N3559, N3558 } = (N114)? { N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231 } : 
                                                                            (N115)? { dcsr_q_xdebugver__31_, dcsr_q_xdebugver__30_, dcsr_q_xdebugver__29_, dcsr_q_xdebugver__28_, dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_, dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_, dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_, dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_, dcsr_q_ebreakm_, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__8_, dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 1'b0;
  assign { N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563 } = (N114)? { N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? dpc_q : 1'b0;
  assign dscratch0_d = (N114)? { N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327 } : 
                       (N115)? dscratch0_q : 1'b0;
  assign dscratch1_d = (N114)? { N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391 } : 
                       (N115)? dscratch1_q : 1'b0;
  assign icache_d = (N114)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423 } : 
                    (N115)? icache_q : 1'b0;
  assign { mstatus_d_sd_, mstatus_d_wpri4__62_, mstatus_d_wpri4__61_, mstatus_d_wpri4__60_, mstatus_d_wpri4__59_, mstatus_d_wpri4__58_, mstatus_d_wpri4__57_, mstatus_d_wpri4__56_, mstatus_d_wpri4__55_, mstatus_d_wpri4__54_, mstatus_d_wpri4__53_, mstatus_d_wpri4__52_, mstatus_d_wpri4__51_, mstatus_d_wpri4__50_, mstatus_d_wpri4__49_, mstatus_d_wpri4__48_, mstatus_d_wpri4__47_, mstatus_d_wpri4__46_, mstatus_d_wpri4__45_, mstatus_d_wpri4__44_, mstatus_d_wpri4__43_, mstatus_d_wpri4__42_, mstatus_d_wpri4__41_, mstatus_d_wpri4__40_, mstatus_d_wpri4__39_, mstatus_d_wpri4__38_, mstatus_d_wpri4__37_, mstatus_d_wpri4__36_, mstatus_d_wpri3__8_, mstatus_d_wpri3__7_, mstatus_d_wpri3__6_, mstatus_d_wpri3__5_, mstatus_d_wpri3__4_, mstatus_d_wpri3__3_, mstatus_d_wpri3__2_, mstatus_d_wpri3__1_, mstatus_d_wpri3__0_, mstatus_d_tsr_, mstatus_d_tw_, mstatus_d_tvm_, mstatus_d_mxr_, mstatus_d_sum_, mstatus_d_mprv_, mstatus_d_xs__1_, mstatus_d_xs__0_, mstatus_d_fs__1_, mstatus_d_fs__0_, N3633, N3632, mstatus_d_wpri2__1_, mstatus_d_wpri2__0_, N3631, N3630, mstatus_d_wpri1_, N3629, mstatus_d_upie_, N3628, mstatus_d_wpri0_, N3627, mstatus_d_uie_ } = (N114)? { N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N115)? { mstatus_q_sd_, mstatus_q_wpri4__62_, mstatus_q_wpri4__61_, mstatus_q_wpri4__60_, mstatus_q_wpri4__59_, mstatus_q_wpri4__58_, mstatus_q_wpri4__57_, mstatus_q_wpri4__56_, mstatus_q_wpri4__55_, mstatus_q_wpri4__54_, mstatus_q_wpri4__53_, mstatus_q_wpri4__52_, mstatus_q_wpri4__51_, mstatus_q_wpri4__50_, mstatus_q_wpri4__49_, mstatus_q_wpri4__48_, mstatus_q_wpri4__47_, mstatus_q_wpri4__46_, mstatus_q_wpri4__45_, mstatus_q_wpri4__44_, mstatus_q_wpri4__43_, mstatus_q_wpri4__42_, mstatus_q_wpri4__41_, mstatus_q_wpri4__40_, mstatus_q_wpri4__39_, mstatus_q_wpri4__38_, mstatus_q_wpri4__37_, mstatus_q_wpri4__36_, mstatus_q_wpri3__8_, mstatus_q_wpri3__7_, mstatus_q_wpri3__6_, mstatus_q_wpri3__5_, mstatus_q_wpri3__4_, mstatus_q_wpri3__3_, mstatus_q_wpri3__2_, mstatus_q_wpri3__1_, mstatus_q_wpri3__0_, tsr_o, tw_o, tvm_o, mxr_o, sum_o, mstatus_q_mprv_, mstatus_q_xs__1_, mstatus_q_xs__0_, fs_o, mstatus_q_mpp__1_, mstatus_q_mpp__0_, mstatus_q_wpri2__1_, mstatus_q_wpri2__0_, mstatus_q_spp_, mstatus_q_mpie_, mstatus_q_wpri1_, mstatus_q_spie_, mstatus_q_upie_, mstatus_q_mie_, mstatus_q_wpri0_, mstatus_q_sie_, mstatus_q_uie_ } : 1'b0;
  assign mie_d = (N114)? { N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515 } : 
                 (N115)? mie_q : 1'b0;
  assign { mip_d_9, mip_d_5, mip_d_1 } = (N114)? { N2581, N2580, N2579 } : 
                                         (N115)? { mip_q_9, mip_q_5, mip_q_1 } : 1'b0;
  assign stvec_d = (N114)? { N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582 } : 
                   (N115)? stvec_q : 1'b0;
  assign sscratch_d = (N114)? { N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646 } : 
                      (N115)? sscratch_q : 1'b0;
  assign { N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634 } = (N114)? { N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? sepc_q : 1'b0;
  assign { N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698 } = (N114)? { N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? scause_q : 1'b0;
  assign { N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762 } = (N114)? { N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? stval_q : 1'b0;
  assign satp_d = (N114)? { N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902 } : 
                  (N115)? { satp_q_mode__3_, satp_q_mode__2_, satp_q_mode__1_, satp_q_mode__0_, satp_q_asid__15_, satp_q_asid__14_, satp_q_asid__13_, satp_q_asid__12_, satp_q_asid__11_, satp_q_asid__10_, satp_q_asid__9_, satp_q_asid__8_, satp_q_asid__7_, satp_q_asid__6_, satp_q_asid__5_, satp_q_asid__4_, satp_q_asid__3_, satp_q_asid__2_, satp_q_asid__1_, asid_o[0:0], satp_ppn_o } : 1'b0;
  assign { medeleg_d[15:15], medeleg_d[13:12], medeleg_d[8:8], medeleg_d[3:3], medeleg_d[0:0] } = (N114)? { N2971, N2970, N2969, N2968, N2967, N2966 } : 
                                                                                                  (N115)? { medeleg_q_15, medeleg_q, medeleg_q_8, medeleg_q_3, medeleg_q_0 } : 1'b0;
  assign { mideleg_d[9:9], mideleg_d[5:5], mideleg_d[1:1] } = (N114)? { N2974, N2973, N2972 } : 
                                                              (N115)? { mideleg_q[9:9], mideleg_q_5, mideleg_q_1 } : 1'b0;
  assign mtvec_d = (N114)? { N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975 } : 
                   (N115)? { N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486 } : 1'b0;
  assign mscratch_d = (N114)? { N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039 } : 
                      (N115)? mscratch_q : 1'b0;
  assign { N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826 } = (N114)? { N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? mepc_q : 1'b0;
  assign { N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890 } = (N114)? { N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? mcause_q : 1'b0;
  assign { N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954 } = (N114)? { N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N115)? mtval_q : 1'b0;
  assign cycle_d = (N114)? { N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295 } : 
                   (N115)? { N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357 } : 1'b0;
  assign dcache_d = (N114)? { N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359 } : 
                    (N115)? { dcache_q, dcache_en_o } : 1'b0;
  assign { fcsr_d_fflags__4_, fcsr_d_fflags__3_, fcsr_d_fflags__2_, fcsr_d_fflags__1_, fcsr_d_fflags__0_ } = (N116)? { N4019, N4020, N4021, N4022, N4023 } : 
                                                                                                             (N117)? { N3557, N3556, N3555, N3554, N3553 } : 1'b0;
  assign N116 = csr_write_fflags_i;
  assign N117 = N4018;
  assign N4160 = (N118)? N5562 : 
                 (N4159)? 1'b1 : 1'b0;
  assign N118 = N4158;
  assign { N4167, N4166, N4165, N4164, N4163, N4162, N4161 } = (N119)? { N3633, N3632, priv_lvl_q[0:0], N3630, mstatus_q_sie_, N3628, 1'b0 } : 
                                                               (N120)? { priv_lvl_q, N3631, mstatus_q_mie_, N3629, 1'b0, N3627 } : 1'b0;
  assign N119 = N5521;
  assign N120 = N4160;
  assign { N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168 } = (N119)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? { N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698 } : 1'b0;
  assign { N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232 } = (N119)? pc_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? { N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634 } : 1'b0;
  assign { N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296 } = (N119)? ex_i[64:1] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? { N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762 } : 1'b0;
  assign { N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360 } = (N119)? { N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? ex_i[128:65] : 1'b0;
  assign { N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424 } = (N119)? { N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? pc_i : 1'b0;
  assign { N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488 } = (N119)? { N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? ex_i[64:1] : 1'b0;
  assign flush_o = (N121)? 1'b0 : 
                   (N4025)? N3552 : 1'b0;
  assign N121 = N4024;
  assign trap_to_priv_lvl[1] = (N121)? N4160 : 
                               (N4025)? 1'b1 : 1'b0;
  assign { N4553, N4552 } = (N121)? { N4160, 1'b1 } : 
                            (N4025)? priv_lvl_q : 1'b0;
  assign mtval_d = (N121)? { N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488 } : 
                   (N4025)? { N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954 } : 1'b0;
  assign { N4560, N4559, N4558, N4557, N4556, N4555, N4554 } = (N121)? { N4167, N4166, N4165, N4164, N4163, N4162, N4161 } : 
                                                               (N4025)? { N3633, N3632, N3631, N3630, N3629, N3628, N3627 } : 1'b0;
  assign scause_d = (N121)? { N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168 } : 
                    (N4025)? { N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698 } : 1'b0;
  assign sepc_d = (N121)? { N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232 } : 
                  (N4025)? { N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634 } : 1'b0;
  assign stval_d = (N121)? { N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296 } : 
                   (N4025)? { N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762 } : 1'b0;
  assign mcause_d = (N121)? { N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360 } : 
                    (N4025)? { N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890 } : 1'b0;
  assign mepc_d = (N121)? { N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424 } : 
                  (N4025)? { N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826 } : 1'b0;
  assign N4571 = (N122)? dcsr_q_ebreakm_ : 
                 (N123)? dcsr_q_ebreaks_ : 
                 (N124)? dcsr_q_ebreaku_ : 
                 (N125)? debug_mode_o : 1'b0;
  assign N122 = N4564;
  assign N123 = N4566;
  assign N124 = N4568;
  assign N125 = N4570;
  assign N4572 = (N122)? dcsr_q_ebreakm_ : 
                 (N123)? dcsr_q_ebreaks_ : 
                 (N124)? dcsr_q_ebreaku_ : 
                 (N125)? 1'b0 : 1'b0;
  assign N4573 = (N126)? N4572 : 
                 (N4563)? 1'b0 : 1'b0;
  assign N126 = N4562;
  assign N4574 = (N126)? N4571 : 
                 (N4563)? debug_mode_o : 1'b0;
  assign { N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575 } = (N126)? pc_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4563)? { N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563 } : 1'b0;
  assign { N4641, N4640, N4639 } = (N126)? { 1'b0, 1'b0, 1'b1 } : 
                                   (N4563)? { N3562, N3561, N3560 } : 1'b0;
  assign { N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644 } = (N127)? pc_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4643)? { N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575 } : 1'b0;
  assign N127 = N4642;
  assign N4708 = (N127)? 1'b1 : 
                 (N4643)? N4574 : 1'b0;
  assign N4709 = (N127)? 1'b1 : 
                 (N4643)? N4573 : 1'b0;
  assign { N4712, N4711, N4710 } = (N127)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N4643)? { N4641, N4640, N4639 } : 1'b0;
  assign N4718 = ~commit_instr_i[0];
  assign { N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783 } = (N128)? commit_instr_i[67:4] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4931)? { trap_vector_base_o[63:2], 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4717)? { N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719 } : 1'b0;
  assign N128 = N5542;
  assign { N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847 } = (N129)? { N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4714)? { N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644 } : 1'b0;
  assign N129 = N4713;
  assign N4911 = (N129)? 1'b1 : 
                 (N4714)? N4708 : 1'b0;
  assign N4912 = (N129)? 1'b1 : 
                 (N4714)? N4709 : 1'b0;
  assign { N4915, N4914, N4913 } = (N129)? { 1'b1, 1'b0, 1'b0 } : 
                                   (N4714)? { N4712, N4711, N4710 } : 1'b0;
  assign { dcsr_d[8:6], dcsr_d[1:0] } = (N60)? { N4915, N4914, N4913, priv_lvl_o } : 
                                        (N61)? { N3562, N3561, N3560, N3559, N3558 } : 1'b0;
  assign dpc_d = (N60)? { N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847 } : 
                 (N61)? { N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563 } : 1'b0;
  assign N4916 = (N60)? N4912 : 
                 (N61)? 1'b0 : 1'b0;
  assign N4917 = (N60)? N4911 : 
                 (N61)? debug_mode_o : 1'b0;
  assign set_debug_pc_o = (N130)? 1'b1 : 
                          (N4919)? N4916 : 1'b0;
  assign N130 = N4918;
  assign en_ld_st_translation_d = (N131)? 1'b1 : 
                                  (N4921)? en_translation_o : 1'b0;
  assign N131 = N4920;
  assign ld_st_priv_lvl_o = (N132)? { mstatus_q_mpp__1_, mstatus_q_mpp__0_ } : 
                            (N133)? priv_lvl_o : 1'b0;
  assign N132 = mprv;
  assign N133 = N4922;
  assign { mstatus_d_mpp__1_, mstatus_d_mpp__0_, mstatus_d_mpie_, mstatus_d_mie_ } = (N134)? { 1'b0, 1'b0, 1'b1, mstatus_q_mpie_ } : 
                                                                                     (N135)? { N4560, N4559, N4557, N4555 } : 1'b0;
  assign N134 = mret;
  assign N135 = N4923;
  assign { N4925, N4924 } = (N134)? { mstatus_q_mpp__1_, mstatus_q_mpp__0_ } : 
                            (N135)? { N4553, N4552 } : 1'b0;
  assign N4927 = (N136)? 1'b1 : 
                 (N137)? mret : 1'b0;
  assign N136 = sret;
  assign N137 = N4926;
  assign { mstatus_d_spp_, mstatus_d_spie_, mstatus_d_sie_ } = (N136)? { 1'b0, 1'b1, mstatus_q_spie_ } : 
                                                               (N137)? { N4558, N4556, N4554 } : 1'b0;
  assign { N4929, N4928 } = (N136)? { 1'b0, mstatus_q_spp_ } : 
                            (N137)? { N4925, N4924 } : 1'b0;
  assign eret_o = (N138)? 1'b1 : 
                  (N139)? N4927 : 1'b0;
  assign N138 = dret;
  assign N139 = N4930;
  assign priv_lvl_d = (N138)? { dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                      (N139)? { N4929, N4928 } : 1'b0;
  assign debug_mode_d = (N138)? 1'b0 : 
                        (N139)? N4917 : 1'b0;
  assign { N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099 } = (N140)? csr_wdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N141)? { N4971, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008, N5009, N5010, N5011, N5012, N5013, N5014, N5015, N5016, N5017, N5018, N5019, N5020, N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028, N5029, N5030, N5031, N5032, N5033, N5034 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N142)? { N5035, N5036, N5037, N5038, N5039, N5040, N5041, N5042, N5043, N5044, N5045, N5046, N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N143)? csr_wdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N144)? csr_wdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N145)? csr_wdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N146)? csr_wdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4970)? csr_wdata_i : 1'b0;
  assign N140 = N4934;
  assign N141 = N4936;
  assign N142 = N4943;
  assign N143 = N4947;
  assign N144 = N4951;
  assign N145 = N4957;
  assign N146 = N4963;
  assign N5163 = (N140)? 1'b1 : 
                 (N141)? 1'b1 : 
                 (N142)? 1'b1 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b0 : 
                 (N4970)? 1'b0 : 1'b0;
  assign N5164 = (N140)? 1'b1 : 
                 (N141)? 1'b1 : 
                 (N142)? 1'b1 : 
                 (N143)? 1'b1 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b0 : 
                 (N4970)? 1'b0 : 1'b0;
  assign N5165 = (N140)? 1'b0 : 
                 (N141)? 1'b0 : 
                 (N142)? 1'b0 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b1 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b0 : 
                 (N4970)? 1'b0 : 1'b0;
  assign N5166 = (N140)? 1'b0 : 
                 (N141)? 1'b0 : 
                 (N142)? 1'b0 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b1 : 
                 (N146)? 1'b0 : 
                 (N4970)? 1'b0 : 1'b0;
  assign N5167 = (N140)? 1'b0 : 
                 (N141)? 1'b0 : 
                 (N142)? 1'b0 : 
                 (N143)? 1'b0 : 
                 (N144)? 1'b0 : 
                 (N145)? 1'b0 : 
                 (N146)? 1'b1 : 
                 (N4970)? 1'b0 : 1'b0;
  assign N5168 = (N147)? N5166 : 
                 (N148)? 1'b0 : 1'b0;
  assign N147 = N4932;
  assign N148 = csr_op_i[6];
  assign N5169 = (N147)? N5167 : 
                 (N148)? 1'b0 : 1'b0;
  assign csr_wdata = (N147)? { N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099 } : 
                     (N148)? csr_wdata_i : 1'b0;
  assign csr_we = (N147)? N5163 : 
                  (N148)? 1'b0 : 1'b0;
  assign csr_read = (N147)? N5164 : 
                    (N148)? 1'b0 : 1'b0;
  assign N5170 = (N147)? N5165 : 
                 (N148)? 1'b0 : 1'b0;
  assign mret = (N149)? 1'b0 : 
                (N5171)? N5168 : 1'b0;
  assign N149 = ex_i[0];
  assign sret = (N149)? 1'b0 : 
                (N5171)? N5170 : 1'b0;
  assign dret = (N149)? 1'b0 : 
                (N5171)? N5169 : 1'b0;
  assign { N5176, N5175 } = (N150)? { 1'b0, 1'b1 } : 
                            (N5174)? { N5172, N5172 } : 1'b0;
  assign N150 = N5173;
  assign { N5180, N5179 } = (N151)? { 1'b0, 1'b1 } : 
                            (N5178)? { N5176, N5175 } : 1'b0;
  assign N151 = N5177;
  assign { N5185, N5184, N5183 } = (N152)? { 1'b0, 1'b1, 1'b1 } : 
                                   (N5182)? { N5177, N5180, N5179 } : 1'b0;
  assign N152 = N5181;
  assign { N5191, N5190, N5189, N5188 } = (N153)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                          (N5187)? { N5185, N5184, N5181, N5183 } : 1'b0;
  assign N153 = N5186;
  assign { N5197, N5196, N5195, N5194 } = (N154)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                          (N5193)? { N5191, N5190, N5189, N5188 } : 1'b0;
  assign N154 = N5192;
  assign N5236 = (N155)? N5235 : 
                 (N5234)? 1'b1 : 1'b0;
  assign N155 = N5233;
  assign { N5241, N5240, N5239, N5238, N5237 } = (N156)? { N5197, N5196, N5195, N5194, N5236 } : 
                                                 (N5200)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N156 = N5199;
  assign { N5252, N5251, N5250, N5249, N5248 } = (N157)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                 (N5247)? { N5241, N5240, N5239, N5238, N5237 } : 1'b0;
  assign N157 = N5246;
  assign { N5259, N5258, N5257, N5256, N5255 } = (N158)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                 (N5254)? { N5252, N5251, N5250, N5249, N5248 } : 1'b0;
  assign N158 = N5253;
  assign { N5264, N5263, N5262, N5261, N5260 } = (N159)? { N5259, N5258, N5257, N5256, N5255 } : 
                                                 (N5243)? { N5241, N5240, N5239, N5238, N5237 } : 1'b0;
  assign N159 = N5242;
  assign { csr_exception_o[128:128], csr_exception_o[68:65], csr_exception_o[0:0] } = (N160)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                                                      (N5266)? { N5261, N5264, N5263, N5262, N5261, N5260 } : 1'b0;
  assign N160 = N5265;
  assign wfi_d = (N161)? 1'b0 : 
                 (N5271)? 1'b1 : 1'b0;
  assign N161 = N5267;
  assign { N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272 } = (N162)? stvec_q[63:2] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N163)? mtvec_q[63:2] : 1'b0;
  assign N162 = N5537;
  assign N163 = trap_to_priv_lvl[1];
  assign { trap_vector_base_o[63:8], N5339, N5338, N5337, N5336, N5335, N5334 } = (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                                  (N60)? { N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272 } : 1'b0;
  assign trap_vector_base_o[7:2] = (N164)? { 1'b0, 1'b0, csr_exception_o[68:65] } : 
                                   (N5341)? { N5339, N5338, N5337, N5336, N5335, N5334 } : 1'b0;
  assign N164 = N5340;
  assign { N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342 } = (N136)? sepc_q : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N137)? mepc_q : 1'b0;
  assign epc_o = (N138)? dpc_q : 
                 (N139)? { N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342 } : 1'b0;
  assign csr_rdata_o[9] = (N165)? N5431 : 
                          (N166)? N5432 : 
                          (N5430)? csr_rdata[9] : 1'b0;
  assign N165 = N5415;
  assign N166 = N5428;
  assign priv_lvl_o = (N61)? { 1'b1, 1'b1 } : 
                      (N60)? priv_lvl_q : 1'b0;
  assign mprv = (N167)? 1'b0 : 
                (N5435)? mstatus_q_mprv_ : 1'b0;
  assign N167 = N5434;
  assign N168 = 1'b0;
  assign N169 = ~csr_read;
  assign N170 = ~csr_addr_i[0];
  assign N179 = ~N178;
  assign N180 = ~csr_addr_i[1];
  assign N188 = ~N187;
  assign N196 = ~N195;
  assign N206 = ~N205;
  assign N215 = ~N214;
  assign N223 = ~N222;
  assign N231 = ~N230;
  assign N239 = ~N238;
  assign N247 = ~N246;
  assign N255 = ~N254;
  assign N263 = ~N262;
  assign N271 = ~N270;
  assign N279 = ~N278;
  assign N280 = ~csr_addr_i[2];
  assign N288 = ~N287;
  assign N296 = ~N295;
  assign N304 = ~N303;
  assign N312 = ~N311;
  assign N320 = ~N319;
  assign N328 = ~N327;
  assign N336 = ~N335;
  assign N344 = ~N343;
  assign N352 = ~N351;
  assign N360 = ~N359;
  assign N368 = ~N367;
  assign N376 = ~N375;
  assign N384 = ~N383;
  assign N392 = ~N391;
  assign N400 = ~N399;
  assign N408 = ~N407;
  assign N416 = ~N415;
  assign N424 = ~N423;
  assign N432 = ~N431;
  assign N440 = ~N439;
  assign N448 = ~N447;
  assign N457 = ~N456;
  assign N465 = ~N464;
  assign N473 = ~N472;
  assign N481 = ~N480;
  assign N490 = ~N489;
  assign N498 = ~N497;
  assign N506 = ~N505;
  assign N514 = ~N513;
  assign N522 = ~N521;
  assign N530 = ~N529;
  assign N566 = ~csr_addr_i[3];
  assign N630 = N5610 | N5611;
  assign N5610 = N5608 | N5609;
  assign N5608 = N5606 | N5607;
  assign N5606 = N5604 | N5605;
  assign N5604 = N5602 | N5603;
  assign N5602 = N5600 | N5601;
  assign N5600 = N5598 | N5599;
  assign N5598 = N5596 | N5597;
  assign N5596 = N5594 | N5595;
  assign N5594 = N5592 | N5593;
  assign N5592 = N5590 | N5591;
  assign N5590 = N5588 | N5589;
  assign N5588 = N5586 | N5587;
  assign N5586 = ~N537;
  assign N5587 = ~N544;
  assign N5589 = ~N551;
  assign N5591 = ~N558;
  assign N5593 = ~N565;
  assign N5595 = ~N573;
  assign N5597 = ~N580;
  assign N5599 = ~N587;
  assign N5601 = ~N594;
  assign N5603 = ~N601;
  assign N5605 = ~N608;
  assign N5607 = ~N615;
  assign N5609 = ~N622;
  assign N5611 = ~N629;
  assign N746 = N631 | N5666;
  assign N5666 = N632 | N5665;
  assign N5665 = N635 | N5664;
  assign N5664 = N637 | N5663;
  assign N5663 = N641 | N5662;
  assign N5662 = N643 | N5661;
  assign N5661 = N645 | N5660;
  assign N5660 = N647 | N5659;
  assign N5659 = N648 | N5658;
  assign N5658 = N649 | N5657;
  assign N5657 = N652 | N5656;
  assign N5656 = N653 | N5655;
  assign N5655 = N656 | N5654;
  assign N5654 = N659 | N5653;
  assign N5653 = N660 | N5652;
  assign N5652 = N661 | N5651;
  assign N5651 = N665 | N5650;
  assign N5650 = N670 | N5649;
  assign N5649 = N675 | N5648;
  assign N5648 = N678 | N5647;
  assign N5647 = N680 | N5646;
  assign N5646 = N681 | N5645;
  assign N5645 = N684 | N5644;
  assign N5644 = N686 | N5643;
  assign N5643 = N687 | N5642;
  assign N5642 = N690 | N5641;
  assign N5641 = N691 | N5640;
  assign N5640 = N692 | N5639;
  assign N5639 = N694 | N5638;
  assign N5638 = N695 | N5637;
  assign N5637 = N696 | N5636;
  assign N5636 = N698 | N5635;
  assign N5635 = N700 | N5634;
  assign N5634 = N701 | N5633;
  assign N5633 = N705 | N5632;
  assign N5632 = N706 | N5631;
  assign N5631 = N707 | N5630;
  assign N5630 = N709 | N5629;
  assign N5629 = N711 | N5628;
  assign N5628 = N714 | N5627;
  assign N5627 = N718 | N5626;
  assign N5626 = N720 | N5625;
  assign N5625 = N723 | N5624;
  assign N5624 = N725 | N5623;
  assign N5623 = N726 | N5622;
  assign N5622 = N728 | N5621;
  assign N5621 = N731 | N5620;
  assign N5620 = N732 | N5619;
  assign N5619 = N734 | N5618;
  assign N5618 = N735 | N5617;
  assign N5617 = N736 | N5616;
  assign N5616 = N737 | N5615;
  assign N5615 = N738 | N5614;
  assign N5614 = N740 | N5613;
  assign N5613 = N741 | N5612;
  assign N5612 = N742 | N745;
  assign N770 = mie_q[63] & mideleg_d[63];
  assign N771 = mie_q[62] & mideleg_d[62];
  assign N772 = mie_q[61] & mideleg_d[61];
  assign N773 = mie_q[60] & mideleg_d[60];
  assign N774 = mie_q[59] & mideleg_d[59];
  assign N775 = mie_q[58] & mideleg_d[58];
  assign N776 = mie_q[57] & mideleg_d[57];
  assign N777 = mie_q[56] & mideleg_d[56];
  assign N778 = mie_q[55] & mideleg_d[55];
  assign N779 = mie_q[54] & mideleg_d[54];
  assign N780 = mie_q[53] & mideleg_d[53];
  assign N781 = mie_q[52] & mideleg_d[52];
  assign N782 = mie_q[51] & mideleg_d[51];
  assign N783 = mie_q[50] & mideleg_d[50];
  assign N784 = mie_q[49] & mideleg_d[49];
  assign N785 = mie_q[48] & mideleg_d[48];
  assign N786 = mie_q[47] & mideleg_d[47];
  assign N787 = mie_q[46] & mideleg_d[46];
  assign N788 = mie_q[45] & mideleg_d[45];
  assign N789 = mie_q[44] & mideleg_d[44];
  assign N790 = mie_q[43] & mideleg_d[43];
  assign N791 = mie_q[42] & mideleg_d[42];
  assign N792 = mie_q[41] & mideleg_d[41];
  assign N793 = mie_q[40] & mideleg_d[40];
  assign N794 = mie_q[39] & mideleg_d[39];
  assign N795 = mie_q[38] & mideleg_d[38];
  assign N796 = mie_q[37] & mideleg_d[37];
  assign N797 = mie_q[36] & mideleg_d[36];
  assign N798 = mie_q[35] & mideleg_d[35];
  assign N799 = mie_q[34] & mideleg_d[34];
  assign N800 = mie_q[33] & mideleg_d[33];
  assign N801 = mie_q[32] & mideleg_d[32];
  assign N802 = mie_q[31] & mideleg_d[31];
  assign N803 = mie_q[30] & mideleg_d[30];
  assign N804 = mie_q[29] & mideleg_d[29];
  assign N805 = mie_q[28] & mideleg_d[28];
  assign N806 = mie_q[27] & mideleg_d[27];
  assign N807 = mie_q[26] & mideleg_d[26];
  assign N808 = mie_q[25] & mideleg_d[25];
  assign N809 = mie_q[24] & mideleg_d[24];
  assign N810 = mie_q[23] & mideleg_d[23];
  assign N811 = mie_q[22] & mideleg_d[22];
  assign N812 = mie_q[21] & mideleg_d[21];
  assign N813 = mie_q[20] & mideleg_d[20];
  assign N814 = mie_q[19] & mideleg_d[19];
  assign N815 = mie_q[18] & mideleg_d[18];
  assign N816 = mie_q[17] & mideleg_d[17];
  assign N817 = mie_q[16] & mideleg_d[16];
  assign N818 = mie_q[15] & mideleg_d[15];
  assign N819 = mie_q[14] & mideleg_d[14];
  assign N820 = mie_q[13] & mideleg_d[13];
  assign N821 = mie_q[12] & mideleg_d[12];
  assign N822 = mie_q[11] & mideleg_d[11];
  assign N823 = mie_q[10] & mideleg_d[10];
  assign N824 = mie_q[9] & mideleg_q[9];
  assign N825 = mie_q[8] & mideleg_d[8];
  assign N826 = mie_q[7] & mideleg_d[7];
  assign N827 = mie_q[6] & mideleg_d[6];
  assign N828 = mie_q[5] & mideleg_q_5;
  assign N829 = mie_q[4] & mideleg_d[4];
  assign N830 = mie_q[3] & mideleg_d[3];
  assign N831 = mie_q[2] & mideleg_d[2];
  assign N832 = mie_q[1] & mideleg_q_1;
  assign N833 = mie_q[0] & mideleg_d[0];
  assign N834 = mip_d[63] & mideleg_d[63];
  assign N835 = mip_d[62] & mideleg_d[62];
  assign N836 = mip_d[61] & mideleg_d[61];
  assign N837 = mip_d[60] & mideleg_d[60];
  assign N838 = mip_d[59] & mideleg_d[59];
  assign N839 = mip_d[58] & mideleg_d[58];
  assign N840 = mip_d[57] & mideleg_d[57];
  assign N841 = mip_d[56] & mideleg_d[56];
  assign N842 = mip_d[55] & mideleg_d[55];
  assign N843 = mip_d[54] & mideleg_d[54];
  assign N844 = mip_d[53] & mideleg_d[53];
  assign N845 = mip_d[52] & mideleg_d[52];
  assign N846 = mip_d[51] & mideleg_d[51];
  assign N847 = mip_d[50] & mideleg_d[50];
  assign N848 = mip_d[49] & mideleg_d[49];
  assign N849 = mip_d[48] & mideleg_d[48];
  assign N850 = mip_d[47] & mideleg_d[47];
  assign N851 = mip_d[46] & mideleg_d[46];
  assign N852 = mip_d[45] & mideleg_d[45];
  assign N853 = mip_d[44] & mideleg_d[44];
  assign N854 = mip_d[43] & mideleg_d[43];
  assign N855 = mip_d[42] & mideleg_d[42];
  assign N856 = mip_d[41] & mideleg_d[41];
  assign N857 = mip_d[40] & mideleg_d[40];
  assign N858 = mip_d[39] & mideleg_d[39];
  assign N859 = mip_d[38] & mideleg_d[38];
  assign N860 = mip_d[37] & mideleg_d[37];
  assign N861 = mip_d[36] & mideleg_d[36];
  assign N862 = mip_d[35] & mideleg_d[35];
  assign N863 = mip_d[34] & mideleg_d[34];
  assign N864 = mip_d[33] & mideleg_d[33];
  assign N865 = mip_d[32] & mideleg_d[32];
  assign N866 = mip_d[31] & mideleg_d[31];
  assign N867 = mip_d[30] & mideleg_d[30];
  assign N868 = mip_d[29] & mideleg_d[29];
  assign N869 = mip_d[28] & mideleg_d[28];
  assign N870 = mip_d[27] & mideleg_d[27];
  assign N871 = mip_d[26] & mideleg_d[26];
  assign N872 = mip_d[25] & mideleg_d[25];
  assign N873 = mip_d[24] & mideleg_d[24];
  assign N874 = mip_d[23] & mideleg_d[23];
  assign N875 = mip_d[22] & mideleg_d[22];
  assign N876 = mip_d[21] & mideleg_d[21];
  assign N877 = mip_d[20] & mideleg_d[20];
  assign N878 = mip_d[19] & mideleg_d[19];
  assign N879 = mip_d[18] & mideleg_d[18];
  assign N880 = mip_d[17] & mideleg_d[17];
  assign N881 = mip_d[16] & mideleg_d[16];
  assign N882 = mip_d[15] & mideleg_d[15];
  assign N883 = mip_d[14] & mideleg_d[14];
  assign N884 = mip_d[13] & mideleg_d[13];
  assign N885 = mip_d[12] & mideleg_d[12];
  assign N886 = mip_q[11] & mideleg_d[11];
  assign N887 = mip_d_10 & mideleg_d[10];
  assign N888 = mip_q_9 & mideleg_q[9];
  assign N889 = mip_d_8 & mideleg_d[8];
  assign N890 = mip_q_7 & mideleg_d[7];
  assign N891 = mip_d_6 & mideleg_d[6];
  assign N892 = mip_q_5 & mideleg_q_5;
  assign N893 = mip_d_4 & mideleg_d[4];
  assign N894 = mip_q_3 & mideleg_d[3];
  assign N895 = mip_d_2 & mideleg_d[2];
  assign N896 = mip_q_1 & mideleg_q_1;
  assign N897 = mip_d_0 & mideleg_d[0];
  assign N898 = N5585 & tvm_o;
  assign N899 = ~N898;
  assign N1029 = ~ex_i[0];
  assign N1030 = ~debug_mode_o;
  assign N1031 = N5667 | N5668;
  assign N5667 = mstatus_q_xs__1_ & mstatus_q_xs__0_;
  assign N5668 = fs_o[1] & fs_o[0];
  assign N1032 = N1030;
  assign N1033 = commit_ack_i[0] & N1029;
  assign N1034 = ~N1033;
  assign N1163 = commit_ack_i[1] & N1029;
  assign N1164 = ~N1163;
  assign N1421 = ~mtvec_rst_load_q;
  assign N1550 = ~csr_we;
  assign N1558 = ~N1557;
  assign N1566 = ~N1565;
  assign N1574 = ~N1573;
  assign N1582 = ~N1581;
  assign N1590 = ~N1589;
  assign N1598 = ~N1597;
  assign N1606 = ~N1605;
  assign N1614 = ~N1613;
  assign N1622 = ~N1621;
  assign N1630 = ~N1629;
  assign N1638 = ~N1637;
  assign N1646 = ~N1645;
  assign N1654 = ~N1653;
  assign N1662 = ~N1661;
  assign N1670 = ~N1669;
  assign N1678 = ~N1677;
  assign N1686 = ~N1685;
  assign N1694 = ~N1693;
  assign N1702 = ~N1701;
  assign N1710 = ~N1709;
  assign N1718 = ~N1717;
  assign N1726 = ~N1725;
  assign N1734 = ~N1733;
  assign N1742 = ~N1741;
  assign N1750 = ~N1749;
  assign N1758 = ~N1757;
  assign N1766 = ~N1765;
  assign N1774 = ~N1773;
  assign N1782 = ~N1781;
  assign N1790 = ~N1789;
  assign N1798 = ~N1797;
  assign N1806 = ~N1805;
  assign N1814 = ~N1813;
  assign N1822 = ~N1821;
  assign N1830 = ~N1829;
  assign N1838 = ~N1837;
  assign N1846 = ~N1845;
  assign N1856 = ~N1855;
  assign N1857 = ~csr_addr_i[11];
  assign N1946 = N5689 | N5690;
  assign N5689 = N5687 | N5688;
  assign N5687 = N5685 | N5686;
  assign N5685 = N5683 | N5684;
  assign N5683 = N5681 | N5682;
  assign N5681 = N5679 | N5680;
  assign N5679 = N5677 | N5678;
  assign N5677 = N5675 | N5676;
  assign N5675 = N5673 | N5674;
  assign N5673 = N5671 | N5672;
  assign N5671 = N5669 | N5670;
  assign N5669 = ~N1868;
  assign N5670 = ~N1875;
  assign N5672 = ~N1882;
  assign N5674 = ~N1889;
  assign N5676 = ~N1896;
  assign N5678 = ~N1903;
  assign N5680 = ~N1910;
  assign N5682 = ~N1917;
  assign N5684 = ~N1924;
  assign N5686 = ~N1931;
  assign N5688 = ~N1938;
  assign N5690 = ~N1945;
  assign N1947 = N1566 | N1558;
  assign N1948 = N1574 | N1947;
  assign N1949 = N1582 | N1948;
  assign N1950 = N1590 | N1949;
  assign N1951 = N1598 | N1950;
  assign N1952 = N1606 | N1951;
  assign N1953 = N1614 | N1952;
  assign N1954 = N1622 | N1953;
  assign N1955 = N1630 | N1954;
  assign N1956 = N1638 | N1955;
  assign N1957 = N1646 | N1956;
  assign N1958 = N1654 | N1957;
  assign N1959 = N1662 | N1958;
  assign N1960 = N1670 | N1959;
  assign N1961 = N1678 | N1960;
  assign N1962 = N1686 | N1961;
  assign N1963 = N1694 | N1962;
  assign N1964 = N1702 | N1963;
  assign N1965 = N1710 | N1964;
  assign N1966 = N1718 | N1965;
  assign N1967 = N1726 | N1966;
  assign N1968 = N1734 | N1967;
  assign N1969 = N1742 | N1968;
  assign N1970 = N1750 | N1969;
  assign N1971 = N1758 | N1970;
  assign N1972 = N1766 | N1971;
  assign N1973 = N1774 | N1972;
  assign N1974 = N1782 | N1973;
  assign N1975 = N1790 | N1974;
  assign N1976 = N1798 | N1975;
  assign N1977 = N1806 | N1976;
  assign N1978 = N1814 | N1977;
  assign N1979 = N1822 | N1978;
  assign N1980 = N1830 | N1979;
  assign N1981 = N1838 | N1980;
  assign N1982 = N1846 | N1981;
  assign N1983 = N1856 | N1982;
  assign N1984 = N1946 | N1983;
  assign N1985 = ~N1984;
  assign N2009 = N5692 | N5693;
  assign N5692 = mie_q[63] & N5691;
  assign N5691 = ~mideleg_d[63];
  assign N5693 = csr_wdata[63] & mideleg_d[63];
  assign N2010 = N5695 | N5696;
  assign N5695 = mie_q[62] & N5694;
  assign N5694 = ~mideleg_d[62];
  assign N5696 = csr_wdata[62] & mideleg_d[62];
  assign N2011 = N5698 | N5699;
  assign N5698 = mie_q[61] & N5697;
  assign N5697 = ~mideleg_d[61];
  assign N5699 = csr_wdata[61] & mideleg_d[61];
  assign N2012 = N5701 | N5702;
  assign N5701 = mie_q[60] & N5700;
  assign N5700 = ~mideleg_d[60];
  assign N5702 = csr_wdata[60] & mideleg_d[60];
  assign N2013 = N5704 | N5705;
  assign N5704 = mie_q[59] & N5703;
  assign N5703 = ~mideleg_d[59];
  assign N5705 = csr_wdata[59] & mideleg_d[59];
  assign N2014 = N5707 | N5708;
  assign N5707 = mie_q[58] & N5706;
  assign N5706 = ~mideleg_d[58];
  assign N5708 = csr_wdata[58] & mideleg_d[58];
  assign N2015 = N5710 | N5711;
  assign N5710 = mie_q[57] & N5709;
  assign N5709 = ~mideleg_d[57];
  assign N5711 = csr_wdata[57] & mideleg_d[57];
  assign N2016 = N5713 | N5714;
  assign N5713 = mie_q[56] & N5712;
  assign N5712 = ~mideleg_d[56];
  assign N5714 = csr_wdata[56] & mideleg_d[56];
  assign N2017 = N5716 | N5717;
  assign N5716 = mie_q[55] & N5715;
  assign N5715 = ~mideleg_d[55];
  assign N5717 = csr_wdata[55] & mideleg_d[55];
  assign N2018 = N5719 | N5720;
  assign N5719 = mie_q[54] & N5718;
  assign N5718 = ~mideleg_d[54];
  assign N5720 = csr_wdata[54] & mideleg_d[54];
  assign N2019 = N5722 | N5723;
  assign N5722 = mie_q[53] & N5721;
  assign N5721 = ~mideleg_d[53];
  assign N5723 = csr_wdata[53] & mideleg_d[53];
  assign N2020 = N5725 | N5726;
  assign N5725 = mie_q[52] & N5724;
  assign N5724 = ~mideleg_d[52];
  assign N5726 = csr_wdata[52] & mideleg_d[52];
  assign N2021 = N5728 | N5729;
  assign N5728 = mie_q[51] & N5727;
  assign N5727 = ~mideleg_d[51];
  assign N5729 = csr_wdata[51] & mideleg_d[51];
  assign N2022 = N5731 | N5732;
  assign N5731 = mie_q[50] & N5730;
  assign N5730 = ~mideleg_d[50];
  assign N5732 = csr_wdata[50] & mideleg_d[50];
  assign N2023 = N5734 | N5735;
  assign N5734 = mie_q[49] & N5733;
  assign N5733 = ~mideleg_d[49];
  assign N5735 = csr_wdata[49] & mideleg_d[49];
  assign N2024 = N5737 | N5738;
  assign N5737 = mie_q[48] & N5736;
  assign N5736 = ~mideleg_d[48];
  assign N5738 = csr_wdata[48] & mideleg_d[48];
  assign N2025 = N5740 | N5741;
  assign N5740 = mie_q[47] & N5739;
  assign N5739 = ~mideleg_d[47];
  assign N5741 = csr_wdata[47] & mideleg_d[47];
  assign N2026 = N5743 | N5744;
  assign N5743 = mie_q[46] & N5742;
  assign N5742 = ~mideleg_d[46];
  assign N5744 = csr_wdata[46] & mideleg_d[46];
  assign N2027 = N5746 | N5747;
  assign N5746 = mie_q[45] & N5745;
  assign N5745 = ~mideleg_d[45];
  assign N5747 = csr_wdata[45] & mideleg_d[45];
  assign N2028 = N5749 | N5750;
  assign N5749 = mie_q[44] & N5748;
  assign N5748 = ~mideleg_d[44];
  assign N5750 = csr_wdata[44] & mideleg_d[44];
  assign N2029 = N5752 | N5753;
  assign N5752 = mie_q[43] & N5751;
  assign N5751 = ~mideleg_d[43];
  assign N5753 = csr_wdata[43] & mideleg_d[43];
  assign N2030 = N5755 | N5756;
  assign N5755 = mie_q[42] & N5754;
  assign N5754 = ~mideleg_d[42];
  assign N5756 = csr_wdata[42] & mideleg_d[42];
  assign N2031 = N5758 | N5759;
  assign N5758 = mie_q[41] & N5757;
  assign N5757 = ~mideleg_d[41];
  assign N5759 = csr_wdata[41] & mideleg_d[41];
  assign N2032 = N5761 | N5762;
  assign N5761 = mie_q[40] & N5760;
  assign N5760 = ~mideleg_d[40];
  assign N5762 = csr_wdata[40] & mideleg_d[40];
  assign N2033 = N5764 | N5765;
  assign N5764 = mie_q[39] & N5763;
  assign N5763 = ~mideleg_d[39];
  assign N5765 = csr_wdata[39] & mideleg_d[39];
  assign N2034 = N5767 | N5768;
  assign N5767 = mie_q[38] & N5766;
  assign N5766 = ~mideleg_d[38];
  assign N5768 = csr_wdata[38] & mideleg_d[38];
  assign N2035 = N5770 | N5771;
  assign N5770 = mie_q[37] & N5769;
  assign N5769 = ~mideleg_d[37];
  assign N5771 = csr_wdata[37] & mideleg_d[37];
  assign N2036 = N5773 | N5774;
  assign N5773 = mie_q[36] & N5772;
  assign N5772 = ~mideleg_d[36];
  assign N5774 = csr_wdata[36] & mideleg_d[36];
  assign N2037 = N5776 | N5777;
  assign N5776 = mie_q[35] & N5775;
  assign N5775 = ~mideleg_d[35];
  assign N5777 = csr_wdata[35] & mideleg_d[35];
  assign N2038 = N5779 | N5780;
  assign N5779 = mie_q[34] & N5778;
  assign N5778 = ~mideleg_d[34];
  assign N5780 = csr_wdata[34] & mideleg_d[34];
  assign N2039 = N5782 | N5783;
  assign N5782 = mie_q[33] & N5781;
  assign N5781 = ~mideleg_d[33];
  assign N5783 = csr_wdata[33] & mideleg_d[33];
  assign N2040 = N5785 | N5786;
  assign N5785 = mie_q[32] & N5784;
  assign N5784 = ~mideleg_d[32];
  assign N5786 = csr_wdata[32] & mideleg_d[32];
  assign N2041 = N5788 | N5789;
  assign N5788 = mie_q[31] & N5787;
  assign N5787 = ~mideleg_d[31];
  assign N5789 = csr_wdata[31] & mideleg_d[31];
  assign N2042 = N5791 | N5792;
  assign N5791 = mie_q[30] & N5790;
  assign N5790 = ~mideleg_d[30];
  assign N5792 = csr_wdata[30] & mideleg_d[30];
  assign N2043 = N5794 | N5795;
  assign N5794 = mie_q[29] & N5793;
  assign N5793 = ~mideleg_d[29];
  assign N5795 = csr_wdata[29] & mideleg_d[29];
  assign N2044 = N5797 | N5798;
  assign N5797 = mie_q[28] & N5796;
  assign N5796 = ~mideleg_d[28];
  assign N5798 = csr_wdata[28] & mideleg_d[28];
  assign N2045 = N5800 | N5801;
  assign N5800 = mie_q[27] & N5799;
  assign N5799 = ~mideleg_d[27];
  assign N5801 = csr_wdata[27] & mideleg_d[27];
  assign N2046 = N5803 | N5804;
  assign N5803 = mie_q[26] & N5802;
  assign N5802 = ~mideleg_d[26];
  assign N5804 = csr_wdata[26] & mideleg_d[26];
  assign N2047 = N5806 | N5807;
  assign N5806 = mie_q[25] & N5805;
  assign N5805 = ~mideleg_d[25];
  assign N5807 = csr_wdata[25] & mideleg_d[25];
  assign N2048 = N5809 | N5810;
  assign N5809 = mie_q[24] & N5808;
  assign N5808 = ~mideleg_d[24];
  assign N5810 = csr_wdata[24] & mideleg_d[24];
  assign N2049 = N5812 | N5813;
  assign N5812 = mie_q[23] & N5811;
  assign N5811 = ~mideleg_d[23];
  assign N5813 = csr_wdata[23] & mideleg_d[23];
  assign N2050 = N5815 | N5816;
  assign N5815 = mie_q[22] & N5814;
  assign N5814 = ~mideleg_d[22];
  assign N5816 = csr_wdata[22] & mideleg_d[22];
  assign N2051 = N5818 | N5819;
  assign N5818 = mie_q[21] & N5817;
  assign N5817 = ~mideleg_d[21];
  assign N5819 = csr_wdata[21] & mideleg_d[21];
  assign N2052 = N5821 | N5822;
  assign N5821 = mie_q[20] & N5820;
  assign N5820 = ~mideleg_d[20];
  assign N5822 = csr_wdata[20] & mideleg_d[20];
  assign N2053 = N5824 | N5825;
  assign N5824 = mie_q[19] & N5823;
  assign N5823 = ~mideleg_d[19];
  assign N5825 = csr_wdata[19] & mideleg_d[19];
  assign N2054 = N5827 | N5828;
  assign N5827 = mie_q[18] & N5826;
  assign N5826 = ~mideleg_d[18];
  assign N5828 = csr_wdata[18] & mideleg_d[18];
  assign N2055 = N5830 | N5831;
  assign N5830 = mie_q[17] & N5829;
  assign N5829 = ~mideleg_d[17];
  assign N5831 = csr_wdata[17] & mideleg_d[17];
  assign N2056 = N5833 | N5834;
  assign N5833 = mie_q[16] & N5832;
  assign N5832 = ~mideleg_d[16];
  assign N5834 = csr_wdata[16] & mideleg_d[16];
  assign N2057 = N5836 | N5837;
  assign N5836 = mie_q[15] & N5835;
  assign N5835 = ~mideleg_d[15];
  assign N5837 = csr_wdata[15] & mideleg_d[15];
  assign N2058 = N5839 | N5840;
  assign N5839 = mie_q[14] & N5838;
  assign N5838 = ~mideleg_d[14];
  assign N5840 = csr_wdata[14] & mideleg_d[14];
  assign N2059 = N5842 | N5843;
  assign N5842 = mie_q[13] & N5841;
  assign N5841 = ~mideleg_d[13];
  assign N5843 = csr_wdata[13] & mideleg_d[13];
  assign N2060 = N5845 | N5846;
  assign N5845 = mie_q[12] & N5844;
  assign N5844 = ~mideleg_d[12];
  assign N5846 = csr_wdata[12] & mideleg_d[12];
  assign N2061 = N5848 | N5849;
  assign N5848 = mie_q[11] & N5847;
  assign N5847 = ~mideleg_d[11];
  assign N5849 = csr_wdata[11] & mideleg_d[11];
  assign N2062 = N5851 | N5852;
  assign N5851 = mie_q[10] & N5850;
  assign N5850 = ~mideleg_d[10];
  assign N5852 = csr_wdata[10] & mideleg_d[10];
  assign N2063 = N5854 | N5855;
  assign N5854 = mie_q[9] & N5853;
  assign N5853 = ~mideleg_q[9];
  assign N5855 = csr_wdata[9] & mideleg_q[9];
  assign N2064 = N5857 | N5858;
  assign N5857 = mie_q[8] & N5856;
  assign N5856 = ~mideleg_d[8];
  assign N5858 = csr_wdata[8] & mideleg_d[8];
  assign N2065 = N5860 | N5861;
  assign N5860 = mie_q[7] & N5859;
  assign N5859 = ~mideleg_d[7];
  assign N5861 = csr_wdata[7] & mideleg_d[7];
  assign N2066 = N5863 | N5864;
  assign N5863 = mie_q[6] & N5862;
  assign N5862 = ~mideleg_d[6];
  assign N5864 = csr_wdata[6] & mideleg_d[6];
  assign N2067 = N5866 | N5867;
  assign N5866 = mie_q[5] & N5865;
  assign N5865 = ~mideleg_q_5;
  assign N5867 = csr_wdata[5] & mideleg_q_5;
  assign N2068 = N5869 | N5870;
  assign N5869 = mie_q[4] & N5868;
  assign N5868 = ~mideleg_d[4];
  assign N5870 = csr_wdata[4] & mideleg_d[4];
  assign N2069 = N5872 | N5873;
  assign N5872 = mie_q[3] & N5871;
  assign N5871 = ~mideleg_d[3];
  assign N5873 = csr_wdata[3] & mideleg_d[3];
  assign N2070 = N5875 | N5876;
  assign N5875 = mie_q[2] & N5874;
  assign N5874 = ~mideleg_d[2];
  assign N5876 = csr_wdata[2] & mideleg_d[2];
  assign N2071 = N5878 | N5879;
  assign N5878 = mie_q[1] & N5877;
  assign N5877 = ~mideleg_q_1;
  assign N5879 = csr_wdata[1] & mideleg_q_1;
  assign N2072 = N5881 | N5882;
  assign N5881 = mie_q[0] & N5880;
  assign N5880 = ~mideleg_d[0];
  assign N5882 = csr_wdata[0] & mideleg_d[0];
  assign N2073 = N5883 | N5884;
  assign N5883 = mip_q_1 & N5877;
  assign N5884 = csr_wdata[1] & mideleg_q_1;
  assign N2074 = N5583 & tvm_o;
  assign N2075 = ~N2074;
  assign N2076 = N5531 | N5536;
  assign N2077 = ~N2076;
  assign N2206 = ~csr_wdata[0];
  assign N2223 = N1581;
  assign N4018 = ~csr_write_fflags_i;
  assign N4019 = csr_wdata_i[4] | fflags_o[4];
  assign N4020 = csr_wdata_i[3] | fflags_o[3];
  assign N4021 = csr_wdata_i[2] | fflags_o[2];
  assign N4022 = csr_wdata_i[1] | fflags_o[1];
  assign N4023 = csr_wdata_i[0] | fflags_o[0];
  assign N4024 = N1030 & ex_i[0];
  assign N4025 = ~N4024;
  assign N4026 = ~ex_i[65];
  assign N4027 = ~ex_i[66];
  assign N4028 = N4026 & N4027;
  assign N4029 = N4026 & ex_i[66];
  assign N4030 = ex_i[65] & N4027;
  assign N4031 = ex_i[65] & ex_i[66];
  assign N4032 = ~ex_i[67];
  assign N4033 = N4028 & N4032;
  assign N4034 = N4028 & ex_i[67];
  assign N4035 = N4030 & N4032;
  assign N4036 = N4030 & ex_i[67];
  assign N4037 = N4029 & N4032;
  assign N4038 = N4029 & ex_i[67];
  assign N4039 = N4031 & N4032;
  assign N4040 = N4031 & ex_i[67];
  assign N4041 = ~ex_i[68];
  assign N4042 = N4033 & N4041;
  assign N4043 = N4033 & ex_i[68];
  assign N4044 = N4035 & N4041;
  assign N4045 = N4035 & ex_i[68];
  assign N4046 = N4037 & N4041;
  assign N4047 = N4037 & ex_i[68];
  assign N4048 = N4039 & N4041;
  assign N4049 = N4039 & ex_i[68];
  assign N4050 = N4034 & N4041;
  assign N4051 = N4034 & ex_i[68];
  assign N4052 = N4036 & N4041;
  assign N4053 = N4036 & ex_i[68];
  assign N4054 = N4038 & N4041;
  assign N4055 = N4038 & ex_i[68];
  assign N4056 = N4040 & N4041;
  assign N4057 = N4040 & ex_i[68];
  assign N4058 = ~ex_i[69];
  assign N4059 = N4042 & N4058;
  assign N4060 = N4042 & ex_i[69];
  assign N4061 = N4044 & N4058;
  assign N4062 = N4044 & ex_i[69];
  assign N4063 = N4046 & N4058;
  assign N4064 = N4046 & ex_i[69];
  assign N4065 = N4048 & N4058;
  assign N4066 = N4048 & ex_i[69];
  assign N4067 = N4050 & N4058;
  assign N4068 = N4050 & ex_i[69];
  assign N4069 = N4052 & N4058;
  assign N4070 = N4052 & ex_i[69];
  assign N4071 = N4054 & N4058;
  assign N4072 = N4054 & ex_i[69];
  assign N4073 = N4056 & N4058;
  assign N4074 = N4056 & ex_i[69];
  assign N4075 = N4043 & N4058;
  assign N4076 = N4043 & ex_i[69];
  assign N4077 = N4045 & N4058;
  assign N4078 = N4045 & ex_i[69];
  assign N4079 = N4047 & N4058;
  assign N4080 = N4047 & ex_i[69];
  assign N4081 = N4049 & N4058;
  assign N4082 = N4049 & ex_i[69];
  assign N4083 = N4051 & N4058;
  assign N4084 = N4051 & ex_i[69];
  assign N4085 = N4053 & N4058;
  assign N4086 = N4053 & ex_i[69];
  assign N4087 = N4055 & N4058;
  assign N4088 = N4055 & ex_i[69];
  assign N4089 = N4057 & N4058;
  assign N4090 = N4057 & ex_i[69];
  assign N4091 = ~ex_i[70];
  assign N4092 = N4059 & N4091;
  assign N4093 = N4059 & ex_i[70];
  assign N4094 = N4061 & N4091;
  assign N4095 = N4061 & ex_i[70];
  assign N4096 = N4063 & N4091;
  assign N4097 = N4063 & ex_i[70];
  assign N4098 = N4065 & N4091;
  assign N4099 = N4065 & ex_i[70];
  assign N4100 = N4067 & N4091;
  assign N4101 = N4067 & ex_i[70];
  assign N4102 = N4069 & N4091;
  assign N4103 = N4069 & ex_i[70];
  assign N4104 = N4071 & N4091;
  assign N4105 = N4071 & ex_i[70];
  assign N4106 = N4073 & N4091;
  assign N4107 = N4073 & ex_i[70];
  assign N4108 = N4075 & N4091;
  assign N4109 = N4075 & ex_i[70];
  assign N4110 = N4077 & N4091;
  assign N4111 = N4077 & ex_i[70];
  assign N4112 = N4079 & N4091;
  assign N4113 = N4079 & ex_i[70];
  assign N4114 = N4081 & N4091;
  assign N4115 = N4081 & ex_i[70];
  assign N4116 = N4083 & N4091;
  assign N4117 = N4083 & ex_i[70];
  assign N4118 = N4085 & N4091;
  assign N4119 = N4085 & ex_i[70];
  assign N4120 = N4087 & N4091;
  assign N4121 = N4087 & ex_i[70];
  assign N4122 = N4089 & N4091;
  assign N4123 = N4089 & ex_i[70];
  assign N4124 = N4060 & N4091;
  assign N4125 = N4060 & ex_i[70];
  assign N4126 = N4062 & N4091;
  assign N4127 = N4062 & ex_i[70];
  assign N4128 = N4064 & N4091;
  assign N4129 = N4064 & ex_i[70];
  assign N4130 = N4066 & N4091;
  assign N4131 = N4066 & ex_i[70];
  assign N4132 = N4068 & N4091;
  assign N4133 = N4068 & ex_i[70];
  assign N4134 = N4070 & N4091;
  assign N4135 = N4070 & ex_i[70];
  assign N4136 = N4072 & N4091;
  assign N4137 = N4072 & ex_i[70];
  assign N4138 = N4074 & N4091;
  assign N4139 = N4074 & ex_i[70];
  assign N4140 = N4076 & N4091;
  assign N4141 = N4076 & ex_i[70];
  assign N4142 = N4078 & N4091;
  assign N4143 = N4078 & ex_i[70];
  assign N4144 = N4080 & N4091;
  assign N4145 = N4080 & ex_i[70];
  assign N4146 = N4082 & N4091;
  assign N4147 = N4082 & ex_i[70];
  assign N4148 = N4084 & N4091;
  assign N4149 = N4084 & ex_i[70];
  assign N4150 = N4086 & N4091;
  assign N4151 = N4086 & ex_i[70];
  assign N4152 = N4088 & N4091;
  assign N4153 = N4088 & ex_i[70];
  assign N4154 = N4090 & N4091;
  assign N4155 = N4090 & ex_i[70];
  assign N4158 = N5885 | N5887;
  assign N5885 = ex_i[128] & N4156;
  assign N5887 = N5886 & N4157;
  assign N5886 = ~ex_i[128];
  assign N4159 = ~N4158;
  assign N4561 = N1030;
  assign N4562 = ex_i[0] & N5503;
  assign N4563 = ~N4562;
  assign N4566 = ~N4565;
  assign N4567 = ~priv_lvl_o[1];
  assign N4570 = ~N4569;
  assign N4642 = debug_req_i & commit_instr_i[201];
  assign N4643 = ~N4642;
  assign N4713 = single_step_o & commit_ack_i[0];
  assign N4714 = ~N4713;
  assign N4715 = N4561 & N4713;
  assign N4716 = ex_i[0] | N5542;
  assign N4717 = ~N4716;
  assign N4918 = N5888 & N5503;
  assign N5888 = debug_mode_o & ex_i[0];
  assign N4919 = ~N4918;
  assign N4920 = N5889 & N5510;
  assign N5889 = mprv & N5508;
  assign N4921 = ~N4920;
  assign N4922 = ~mprv;
  assign N4923 = ~mret;
  assign N4926 = ~sret;
  assign N4930 = ~dret;
  assign N4931 = ex_i[0] & N5541;
  assign N4932 = ~csr_op_i[6];
  assign N4934 = ~N4933;
  assign N4936 = ~N4935;
  assign N4937 = ~csr_op_i[5];
  assign N4943 = ~N4942;
  assign N4947 = ~N4946;
  assign N4948 = ~csr_op_i[0];
  assign N4951 = ~N4950;
  assign N4952 = ~csr_op_i[2];
  assign N4957 = ~N4956;
  assign N4963 = ~N4962;
  assign N4964 = N4936 | N4934;
  assign N4965 = N4943 | N4964;
  assign N4966 = N4947 | N4965;
  assign N4967 = N4951 | N4966;
  assign N4968 = N4957 | N4967;
  assign N4969 = N4963 | N4968;
  assign N4970 = ~N4969;
  assign N4971 = csr_wdata_i[63] | csr_rdata_o[63];
  assign N4972 = csr_wdata_i[62] | csr_rdata_o[62];
  assign N4973 = csr_wdata_i[61] | csr_rdata_o[61];
  assign N4974 = csr_wdata_i[60] | csr_rdata_o[60];
  assign N4975 = csr_wdata_i[59] | csr_rdata_o[59];
  assign N4976 = csr_wdata_i[58] | csr_rdata_o[58];
  assign N4977 = csr_wdata_i[57] | csr_rdata_o[57];
  assign N4978 = csr_wdata_i[56] | csr_rdata_o[56];
  assign N4979 = csr_wdata_i[55] | csr_rdata_o[55];
  assign N4980 = csr_wdata_i[54] | csr_rdata_o[54];
  assign N4981 = csr_wdata_i[53] | csr_rdata_o[53];
  assign N4982 = csr_wdata_i[52] | csr_rdata_o[52];
  assign N4983 = csr_wdata_i[51] | csr_rdata_o[51];
  assign N4984 = csr_wdata_i[50] | csr_rdata_o[50];
  assign N4985 = csr_wdata_i[49] | csr_rdata_o[49];
  assign N4986 = csr_wdata_i[48] | csr_rdata_o[48];
  assign N4987 = csr_wdata_i[47] | csr_rdata_o[47];
  assign N4988 = csr_wdata_i[46] | csr_rdata_o[46];
  assign N4989 = csr_wdata_i[45] | csr_rdata_o[45];
  assign N4990 = csr_wdata_i[44] | csr_rdata_o[44];
  assign N4991 = csr_wdata_i[43] | csr_rdata_o[43];
  assign N4992 = csr_wdata_i[42] | csr_rdata_o[42];
  assign N4993 = csr_wdata_i[41] | csr_rdata_o[41];
  assign N4994 = csr_wdata_i[40] | csr_rdata_o[40];
  assign N4995 = csr_wdata_i[39] | csr_rdata_o[39];
  assign N4996 = csr_wdata_i[38] | csr_rdata_o[38];
  assign N4997 = csr_wdata_i[37] | csr_rdata_o[37];
  assign N4998 = csr_wdata_i[36] | csr_rdata_o[36];
  assign N4999 = csr_wdata_i[35] | csr_rdata_o[35];
  assign N5000 = csr_wdata_i[34] | csr_rdata_o[34];
  assign N5001 = csr_wdata_i[33] | csr_rdata_o[33];
  assign N5002 = csr_wdata_i[32] | csr_rdata_o[32];
  assign N5003 = csr_wdata_i[31] | csr_rdata_o[31];
  assign N5004 = csr_wdata_i[30] | csr_rdata_o[30];
  assign N5005 = csr_wdata_i[29] | csr_rdata_o[29];
  assign N5006 = csr_wdata_i[28] | csr_rdata_o[28];
  assign N5007 = csr_wdata_i[27] | csr_rdata_o[27];
  assign N5008 = csr_wdata_i[26] | csr_rdata_o[26];
  assign N5009 = csr_wdata_i[25] | csr_rdata_o[25];
  assign N5010 = csr_wdata_i[24] | csr_rdata_o[24];
  assign N5011 = csr_wdata_i[23] | csr_rdata_o[23];
  assign N5012 = csr_wdata_i[22] | csr_rdata_o[22];
  assign N5013 = csr_wdata_i[21] | csr_rdata_o[21];
  assign N5014 = csr_wdata_i[20] | csr_rdata_o[20];
  assign N5015 = csr_wdata_i[19] | csr_rdata_o[19];
  assign N5016 = csr_wdata_i[18] | csr_rdata_o[18];
  assign N5017 = csr_wdata_i[17] | csr_rdata_o[17];
  assign N5018 = csr_wdata_i[16] | csr_rdata_o[16];
  assign N5019 = csr_wdata_i[15] | csr_rdata_o[15];
  assign N5020 = csr_wdata_i[14] | csr_rdata_o[14];
  assign N5021 = csr_wdata_i[13] | csr_rdata_o[13];
  assign N5022 = csr_wdata_i[12] | csr_rdata_o[12];
  assign N5023 = csr_wdata_i[11] | csr_rdata_o[11];
  assign N5024 = csr_wdata_i[10] | csr_rdata_o[10];
  assign N5025 = csr_wdata_i[9] | csr_rdata[9];
  assign N5026 = csr_wdata_i[8] | csr_rdata_o[8];
  assign N5027 = csr_wdata_i[7] | csr_rdata_o[7];
  assign N5028 = csr_wdata_i[6] | csr_rdata_o[6];
  assign N5029 = csr_wdata_i[5] | csr_rdata_o[5];
  assign N5030 = csr_wdata_i[4] | csr_rdata_o[4];
  assign N5031 = csr_wdata_i[3] | csr_rdata_o[3];
  assign N5032 = csr_wdata_i[2] | csr_rdata_o[2];
  assign N5033 = csr_wdata_i[1] | csr_rdata_o[1];
  assign N5034 = csr_wdata_i[0] | csr_rdata_o[0];
  assign N5035 = N5890 & csr_rdata_o[63];
  assign N5890 = ~csr_wdata_i[63];
  assign N5036 = N5891 & csr_rdata_o[62];
  assign N5891 = ~csr_wdata_i[62];
  assign N5037 = N5892 & csr_rdata_o[61];
  assign N5892 = ~csr_wdata_i[61];
  assign N5038 = N5893 & csr_rdata_o[60];
  assign N5893 = ~csr_wdata_i[60];
  assign N5039 = N5894 & csr_rdata_o[59];
  assign N5894 = ~csr_wdata_i[59];
  assign N5040 = N5895 & csr_rdata_o[58];
  assign N5895 = ~csr_wdata_i[58];
  assign N5041 = N5896 & csr_rdata_o[57];
  assign N5896 = ~csr_wdata_i[57];
  assign N5042 = N5897 & csr_rdata_o[56];
  assign N5897 = ~csr_wdata_i[56];
  assign N5043 = N5898 & csr_rdata_o[55];
  assign N5898 = ~csr_wdata_i[55];
  assign N5044 = N5899 & csr_rdata_o[54];
  assign N5899 = ~csr_wdata_i[54];
  assign N5045 = N5900 & csr_rdata_o[53];
  assign N5900 = ~csr_wdata_i[53];
  assign N5046 = N5901 & csr_rdata_o[52];
  assign N5901 = ~csr_wdata_i[52];
  assign N5047 = N5902 & csr_rdata_o[51];
  assign N5902 = ~csr_wdata_i[51];
  assign N5048 = N5903 & csr_rdata_o[50];
  assign N5903 = ~csr_wdata_i[50];
  assign N5049 = N5904 & csr_rdata_o[49];
  assign N5904 = ~csr_wdata_i[49];
  assign N5050 = N5905 & csr_rdata_o[48];
  assign N5905 = ~csr_wdata_i[48];
  assign N5051 = N5906 & csr_rdata_o[47];
  assign N5906 = ~csr_wdata_i[47];
  assign N5052 = N5907 & csr_rdata_o[46];
  assign N5907 = ~csr_wdata_i[46];
  assign N5053 = N5908 & csr_rdata_o[45];
  assign N5908 = ~csr_wdata_i[45];
  assign N5054 = N5909 & csr_rdata_o[44];
  assign N5909 = ~csr_wdata_i[44];
  assign N5055 = N5910 & csr_rdata_o[43];
  assign N5910 = ~csr_wdata_i[43];
  assign N5056 = N5911 & csr_rdata_o[42];
  assign N5911 = ~csr_wdata_i[42];
  assign N5057 = N5912 & csr_rdata_o[41];
  assign N5912 = ~csr_wdata_i[41];
  assign N5058 = N5913 & csr_rdata_o[40];
  assign N5913 = ~csr_wdata_i[40];
  assign N5059 = N5914 & csr_rdata_o[39];
  assign N5914 = ~csr_wdata_i[39];
  assign N5060 = N5915 & csr_rdata_o[38];
  assign N5915 = ~csr_wdata_i[38];
  assign N5061 = N5916 & csr_rdata_o[37];
  assign N5916 = ~csr_wdata_i[37];
  assign N5062 = N5917 & csr_rdata_o[36];
  assign N5917 = ~csr_wdata_i[36];
  assign N5063 = N5918 & csr_rdata_o[35];
  assign N5918 = ~csr_wdata_i[35];
  assign N5064 = N5919 & csr_rdata_o[34];
  assign N5919 = ~csr_wdata_i[34];
  assign N5065 = N5920 & csr_rdata_o[33];
  assign N5920 = ~csr_wdata_i[33];
  assign N5066 = N5921 & csr_rdata_o[32];
  assign N5921 = ~csr_wdata_i[32];
  assign N5067 = N5922 & csr_rdata_o[31];
  assign N5922 = ~csr_wdata_i[31];
  assign N5068 = N5923 & csr_rdata_o[30];
  assign N5923 = ~csr_wdata_i[30];
  assign N5069 = N5924 & csr_rdata_o[29];
  assign N5924 = ~csr_wdata_i[29];
  assign N5070 = N5925 & csr_rdata_o[28];
  assign N5925 = ~csr_wdata_i[28];
  assign N5071 = N5926 & csr_rdata_o[27];
  assign N5926 = ~csr_wdata_i[27];
  assign N5072 = N5927 & csr_rdata_o[26];
  assign N5927 = ~csr_wdata_i[26];
  assign N5073 = N5928 & csr_rdata_o[25];
  assign N5928 = ~csr_wdata_i[25];
  assign N5074 = N5929 & csr_rdata_o[24];
  assign N5929 = ~csr_wdata_i[24];
  assign N5075 = N5930 & csr_rdata_o[23];
  assign N5930 = ~csr_wdata_i[23];
  assign N5076 = N5931 & csr_rdata_o[22];
  assign N5931 = ~csr_wdata_i[22];
  assign N5077 = N5932 & csr_rdata_o[21];
  assign N5932 = ~csr_wdata_i[21];
  assign N5078 = N5933 & csr_rdata_o[20];
  assign N5933 = ~csr_wdata_i[20];
  assign N5079 = N5934 & csr_rdata_o[19];
  assign N5934 = ~csr_wdata_i[19];
  assign N5080 = N5935 & csr_rdata_o[18];
  assign N5935 = ~csr_wdata_i[18];
  assign N5081 = N5936 & csr_rdata_o[17];
  assign N5936 = ~csr_wdata_i[17];
  assign N5082 = N5937 & csr_rdata_o[16];
  assign N5937 = ~csr_wdata_i[16];
  assign N5083 = N5938 & csr_rdata_o[15];
  assign N5938 = ~csr_wdata_i[15];
  assign N5084 = N5939 & csr_rdata_o[14];
  assign N5939 = ~csr_wdata_i[14];
  assign N5085 = N5940 & csr_rdata_o[13];
  assign N5940 = ~csr_wdata_i[13];
  assign N5086 = N5941 & csr_rdata_o[12];
  assign N5941 = ~csr_wdata_i[12];
  assign N5087 = N5942 & csr_rdata_o[11];
  assign N5942 = ~csr_wdata_i[11];
  assign N5088 = N5943 & csr_rdata_o[10];
  assign N5943 = ~csr_wdata_i[10];
  assign N5089 = N5944 & csr_rdata[9];
  assign N5944 = ~csr_wdata_i[9];
  assign N5090 = N5945 & csr_rdata_o[8];
  assign N5945 = ~csr_wdata_i[8];
  assign N5091 = N5946 & csr_rdata_o[7];
  assign N5946 = ~csr_wdata_i[7];
  assign N5092 = N5947 & csr_rdata_o[6];
  assign N5947 = ~csr_wdata_i[6];
  assign N5093 = N5948 & csr_rdata_o[5];
  assign N5948 = ~csr_wdata_i[5];
  assign N5094 = N5949 & csr_rdata_o[4];
  assign N5949 = ~csr_wdata_i[4];
  assign N5095 = N5950 & csr_rdata_o[3];
  assign N5950 = ~csr_wdata_i[3];
  assign N5096 = N5951 & csr_rdata_o[2];
  assign N5951 = ~csr_wdata_i[2];
  assign N5097 = N5952 & csr_rdata_o[1];
  assign N5952 = ~csr_wdata_i[1];
  assign N5098 = N5953 & csr_rdata_o[0];
  assign N5953 = ~csr_wdata_i[0];
  assign N5171 = ~ex_i[0];
  assign N5172 = mie_q[5] & mip_q_5;
  assign N5173 = mie_q[1] & mip_q_1;
  assign N5174 = ~N5173;
  assign N5177 = mie_q[9] & N5954;
  assign N5954 = mip_q_9 | irq_i[1];
  assign N5178 = ~N5177;
  assign N5181 = mip_q_7 & mie_q[7];
  assign N5182 = ~N5181;
  assign N5186 = mip_q_3 & mie_q[3];
  assign N5187 = ~N5186;
  assign N5192 = mip_q[11] & mie_q[11];
  assign N5193 = ~N5192;
  assign N5198 = N5957 & N5959;
  assign N5957 = N1030 & N5956;
  assign N5956 = N5955 | dcsr_q_stepie_;
  assign N5955 = ~single_step_o;
  assign N5959 = N5958 | N5565;
  assign N5958 = mstatus_q_mie_ & N5563;
  assign N5199 = N5194 & N5198;
  assign N5200 = ~N5199;
  assign N5201 = ~N5194;
  assign N5202 = ~N5195;
  assign N5203 = N5201 & N5202;
  assign N5204 = N5201 & N5195;
  assign N5205 = N5194 & N5202;
  assign N5206 = N5194 & N5195;
  assign N5207 = ~N5196;
  assign N5208 = N5203 & N5207;
  assign N5209 = N5203 & N5196;
  assign N5210 = N5205 & N5207;
  assign N5211 = N5205 & N5196;
  assign N5212 = N5204 & N5207;
  assign N5213 = N5204 & N5196;
  assign N5214 = N5206 & N5207;
  assign N5215 = N5206 & N5196;
  assign N5216 = ~N5197;
  assign N5217 = N5208 & N5216;
  assign N5218 = N5208 & N5197;
  assign N5219 = N5210 & N5216;
  assign N5220 = N5210 & N5197;
  assign N5221 = N5212 & N5216;
  assign N5222 = N5212 & N5197;
  assign N5223 = N5214 & N5216;
  assign N5224 = N5214 & N5197;
  assign N5225 = N5209 & N5216;
  assign N5226 = N5209 & N5197;
  assign N5227 = N5211 & N5216;
  assign N5228 = N5211 & N5197;
  assign N5229 = N5213 & N5216;
  assign N5230 = N5213 & N5197;
  assign N5231 = N5215 & N5216;
  assign N5232 = N5215 & N5197;
  assign N5234 = ~N5233;
  assign N5235 = N5960 | N5547;
  assign N5960 = mstatus_q_sie_ & N5545;
  assign N5242 = csr_we | csr_read;
  assign N5243 = ~N5242;
  assign N5244 = priv_lvl_o[1] & csr_addr_i[9];
  assign N5245 = priv_lvl_o[0] & csr_addr_i[8];
  assign N5247 = ~N5246;
  assign N5253 = N5561 & N1030;
  assign N5254 = ~N5253;
  assign N5265 = update_access_exception | read_access_exception;
  assign N5266 = ~N5265;
  assign N5267 = N6024 | irq_i[1];
  assign N6024 = N6023 | debug_req_i;
  assign N6023 = N6022 | mip_d_0;
  assign N6022 = N6021 | mip_q_1;
  assign N6021 = N6020 | mip_d_2;
  assign N6020 = N6019 | mip_q_3;
  assign N6019 = N6018 | mip_d_4;
  assign N6018 = N6017 | mip_q_5;
  assign N6017 = N6016 | mip_d_6;
  assign N6016 = N6015 | mip_q_7;
  assign N6015 = N6014 | mip_d_8;
  assign N6014 = N6013 | mip_q_9;
  assign N6013 = N6012 | mip_d_10;
  assign N6012 = N6011 | mip_q[11];
  assign N6011 = N6010 | mip_d[12];
  assign N6010 = N6009 | mip_d[13];
  assign N6009 = N6008 | mip_d[14];
  assign N6008 = N6007 | mip_d[15];
  assign N6007 = N6006 | mip_d[16];
  assign N6006 = N6005 | mip_d[17];
  assign N6005 = N6004 | mip_d[18];
  assign N6004 = N6003 | mip_d[19];
  assign N6003 = N6002 | mip_d[20];
  assign N6002 = N6001 | mip_d[21];
  assign N6001 = N6000 | mip_d[22];
  assign N6000 = N5999 | mip_d[23];
  assign N5999 = N5998 | mip_d[24];
  assign N5998 = N5997 | mip_d[25];
  assign N5997 = N5996 | mip_d[26];
  assign N5996 = N5995 | mip_d[27];
  assign N5995 = N5994 | mip_d[28];
  assign N5994 = N5993 | mip_d[29];
  assign N5993 = N5992 | mip_d[30];
  assign N5992 = N5991 | mip_d[31];
  assign N5991 = N5990 | mip_d[32];
  assign N5990 = N5989 | mip_d[33];
  assign N5989 = N5988 | mip_d[34];
  assign N5988 = N5987 | mip_d[35];
  assign N5987 = N5986 | mip_d[36];
  assign N5986 = N5985 | mip_d[37];
  assign N5985 = N5984 | mip_d[38];
  assign N5984 = N5983 | mip_d[39];
  assign N5983 = N5982 | mip_d[40];
  assign N5982 = N5981 | mip_d[41];
  assign N5981 = N5980 | mip_d[42];
  assign N5980 = N5979 | mip_d[43];
  assign N5979 = N5978 | mip_d[44];
  assign N5978 = N5977 | mip_d[45];
  assign N5977 = N5976 | mip_d[46];
  assign N5976 = N5975 | mip_d[47];
  assign N5975 = N5974 | mip_d[48];
  assign N5974 = N5973 | mip_d[49];
  assign N5973 = N5972 | mip_d[50];
  assign N5972 = N5971 | mip_d[51];
  assign N5971 = N5970 | mip_d[52];
  assign N5970 = N5969 | mip_d[53];
  assign N5969 = N5968 | mip_d[54];
  assign N5968 = N5967 | mip_d[55];
  assign N5967 = N5966 | mip_d[56];
  assign N5966 = N5965 | mip_d[57];
  assign N5965 = N5964 | mip_d[58];
  assign N5964 = N5963 | mip_d[59];
  assign N5963 = N5962 | mip_d[60];
  assign N5962 = N5961 | mip_d[61];
  assign N5961 = mip_d[63] | mip_d[62];
  assign N5268 = N6025 & N1029;
  assign N6025 = N1030 & N5520;
  assign N5269 = N5268 | N5267;
  assign N5270 = ~N5267;
  assign N5271 = N5268 & N5270;
  assign N5340 = N6026 & csr_exception_o[128];
  assign N6026 = mtvec_q[0] | stvec_q[0];
  assign N5341 = ~N5340;
  assign N5415 = ~N5414;
  assign N5416 = ~csr_addr_i[6];
  assign N5428 = ~N5427;
  assign N5429 = N5428 | N5415;
  assign N5430 = ~N5429;
  assign N5431 = csr_rdata[9] | irq_i[1];
  assign N5432 = csr_rdata[9] | N6027;
  assign N6027 = irq_i[1] & mideleg_q[9];
  assign N5433 = N5525 & N5527;
  assign en_translation_o = N5433;
  assign icache_en_o = icache_q[0] & N1030;
  assign N5434 = debug_mode_o & N6028;
  assign N6028 = ~dcsr_q_mprven_;
  assign N5435 = ~N5434;
  assign N5436 = ~rst_ni;
  assign N5437 = ~debug_mode_o;

endmodule