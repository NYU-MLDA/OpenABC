module bsg_mem_1r1w_synth_width_p128_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [127:0] w_data_i;
  input [0:0] r_addr_i;
  output [127:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [127:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10;
  wire [255:0] mem;
  reg mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,
  mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,mem_247_sv2v_reg,
  mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,
  mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,
  mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,
  mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,
  mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,
  mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,
  mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,mem_214_sv2v_reg,
  mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,
  mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,
  mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,
  mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,
  mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,
  mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,
  mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,
  mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,
  mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,
  mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,mem_167_sv2v_reg,
  mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,
  mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,
  mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,
  mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,
  mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,
  mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,
  mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,mem_134_sv2v_reg,
  mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,
  mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,
  mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,
  mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,
  mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,
  mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,
  mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,
  mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,
  mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,
  mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,
  mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,
  mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,
  mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,
  mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,
  mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,
  mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,
  mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,
  mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,
  mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,
  mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,
  mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,
  mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,
  mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,
  mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,
  mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,
  mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,
  mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,
  mem_0_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[255] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[254] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[253] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[252] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[251] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[250] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[249] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[248] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[247] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[246] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[245] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[244] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[243] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[242] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[241] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[240] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[239] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[238] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[237] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[236] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[235] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[234] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[233] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[232] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[231] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[230] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[229] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[228] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[227] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[226] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[225] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[224] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[223] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[222] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[221] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[220] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[219] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[218] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[217] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[216] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[215] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[214] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[213] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[212] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[211] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[210] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[209] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[208] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[207] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[206] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[205] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[204] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[203] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[202] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[201] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[200] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[199] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[198] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[197] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[140] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[139] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[138] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[137] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[136] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[135] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[134] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[133] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[132] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[131] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[130] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[129] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[128] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_255_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_254_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_253_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_252_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_251_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_250_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_249_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_248_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_247_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_246_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_245_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_244_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_243_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_242_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_241_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_240_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_239_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_238_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_237_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_236_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_235_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_234_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_233_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_232_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_231_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_230_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_229_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_228_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_227_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_226_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_225_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_224_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_223_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_222_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_221_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_220_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_219_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_218_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_217_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_216_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_215_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_214_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_213_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_212_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_211_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_210_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_209_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_208_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_207_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_206_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_205_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_204_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_203_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_202_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_201_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_200_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_199_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_198_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_197_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_196_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_195_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_194_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_193_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_192_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_191_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_190_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_189_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_188_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_187_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_186_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_185_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_184_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_183_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_182_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_181_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_180_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_179_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_178_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_177_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_176_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_175_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_174_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_173_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_172_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_171_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_170_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_169_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_168_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_167_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_166_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_165_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_164_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_163_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_162_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_161_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_160_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_159_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_158_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_157_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_156_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_155_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_154_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_153_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_152_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_151_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_150_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_149_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_148_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_147_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_146_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_145_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_144_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_143_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_142_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_141_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_140_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_139_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_138_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_137_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_136_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_135_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_134_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_133_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_132_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_131_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_130_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_129_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_128_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_127_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_126_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_125_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_124_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_123_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_122_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_121_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_120_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_119_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_118_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_117_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_116_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_115_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_114_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_113_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_112_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_111_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_110_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_109_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_108_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_107_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_106_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_105_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_104_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_103_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_102_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_101_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_100_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_99_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_98_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_97_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_96_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_95_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_94_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_93_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_92_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_91_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_90_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_89_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_88_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_87_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_86_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_85_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_84_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_83_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_82_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_81_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_80_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_79_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_78_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_77_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_76_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_75_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_74_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_73_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_72_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_71_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_70_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_69_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_68_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_67_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_66_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_65_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_64_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_63_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_62_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N5 = ~w_addr_i[0];
  assign { N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], N5, N5 } : 
                               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

endmodule